module bfloat16_spi_top (clk,
    miso,
    mosi,
    rst,
    ss,
    VPWR,
    VGND);
 input clk;
 output miso;
 input mosi;
 input rst;
 input ss;
 inout VPWR;
 inout VGND;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire net1821;
 wire _01492_;
 wire net1816;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire net74;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_44_clk;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire net64;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire net1775;
 wire _01762_;
 wire _01763_;
 wire net1760;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire net48;
 wire net46;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire net1709;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_7_clk;
 wire _01843_;
 wire _01844_;
 wire clknet_leaf_42_clk;
 wire _01846_;
 wire _01847_;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_36_clk;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire net1691;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_82_clk;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire clknet_leaf_54_clk;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire clknet_leaf_95_clk;
 wire _01946_;
 wire net45;
 wire _01948_;
 wire _01949_;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_93_clk;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_85_clk;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire clknet_leaf_84_clk;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire net1653;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire clknet_leaf_87_clk;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire clknet_leaf_88_clk;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire net1776;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire clknet_leaf_96_clk;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire net50;
 wire net1788;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire net121;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire clknet_leaf_12_clk;
 wire _02248_;
 wire net1703;
 wire _02250_;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_14_clk;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire net1719;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire net1818;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire clknet_leaf_74_clk;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire net1664;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire clknet_leaf_57_clk;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire net1663;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire clknet_leaf_59_clk;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire clknet_leaf_97_clk;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire clknet_leaf_56_clk;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire net49;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire clknet_leaf_61_clk;
 wire _02380_;
 wire _02381_;
 wire clknet_leaf_90_clk;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire net1657;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire net1661;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire clknet_leaf_98_clk;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire net76;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire net1736;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire net1716;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire net1737;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire net75;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire net78;
 wire _02650_;
 wire net1731;
 wire _02652_;
 wire net124;
 wire _02654_;
 wire net1725;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire net123;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_91_clk;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire net1851;
 wire _02726_;
 wire net79;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire clknet_leaf_38_clk;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire net1756;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire net93;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire net1724;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire net1763;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire clknet_leaf_9_clk;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire net1745;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire net1767;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire net1708;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire net1749;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire net1704;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire clknet_leaf_10_clk;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire net129;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire net1715;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire net1793;
 wire _03361_;
 wire net1792;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire net81;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire net1761;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire clknet_leaf_30_clk;
 wire net1683;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire net1755;
 wire _03627_;
 wire _03628_;
 wire net1707;
 wire _03630_;
 wire _03631_;
 wire net94;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire net1759;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire net82;
 wire _03654_;
 wire _03655_;
 wire net65;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire net1689;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire net1671;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire net1649;
 wire _03785_;
 wire net51;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire net1672;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire net1790;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire clknet_leaf_3_clk;
 wire net1754;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire net1698;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire clknet_leaf_31_clk;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire net52;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire net56;
 wire net1772;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire net125;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire clknet_leaf_17_clk;
 wire _04054_;
 wire clknet_leaf_4_clk;
 wire _04056_;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_18_clk;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire net67;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire clknet_leaf_50_clk;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire clknet_leaf_75_clk;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire net1876;
 wire _04130_;
 wire _04131_;
 wire clknet_leaf_47_clk;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire clknet_leaf_76_clk;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire clknet_leaf_99_clk;
 wire _04152_;
 wire net55;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire clknet_leaf_77_clk;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire net1670;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire clknet_leaf_78_clk;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire clknet_leaf_79_clk;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire clknet_leaf_80_clk;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire net68;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire clknet_leaf_100_clk;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire net1824;
 wire _04386_;
 wire net84;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire clknet_leaf_33_clk;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire net1744;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire net1752;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire net1713;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire net95;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire net1750;
 wire _04670_;
 wire net1692;
 wire _04672_;
 wire net1753;
 wire _04674_;
 wire _04675_;
 wire net69;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire net85;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire net1694;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire net1674;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire net117;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire net1764;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire net130;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire net59;
 wire net58;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire net1722;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire net57;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire net133;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire net132;
 wire _05052_;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_21_clk;
 wire _05055_;
 wire clknet_leaf_20_clk;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire net134;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire clknet_leaf_49_clk;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire clknet_leaf_62_clk;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire clknet_leaf_67_clk;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire clknet_leaf_69_clk;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire clknet_leaf_51_clk;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire clknet_leaf_101_clk;
 wire clknet_leaf_66_clk;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire clknet_leaf_68_clk;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire clknet_leaf_70_clk;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire net1658;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire clknet_leaf_71_clk;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire clknet_leaf_102_clk;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire net70;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire net86;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire net96;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire net118;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire net97;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire clknet_leaf_5_clk;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire net71;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire net1769;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire net1665;
 wire _05572_;
 wire _05573_;
 wire net1774;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire net100;
 wire net99;
 wire _05586_;
 wire _05587_;
 wire net1701;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire net126;
 wire _05598_;
 wire _05599_;
 wire clknet_leaf_11_clk;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire net135;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire net136;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire clknet_leaf_39_clk;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire clknet_leaf_52_clk;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire clknet_leaf_72_clk;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire net119;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire clknet_leaf_34_clk;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire net89;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire net88;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire net72;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire net1743;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire net137;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire net91;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire net1739;
 wire _06573_;
 wire _06574_;
 wire net110;
 wire net109;
 wire _06577_;
 wire net127;
 wire net1741;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire net90;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire _06602_;
 wire _06603_;
 wire _06604_;
 wire _06605_;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire _06621_;
 wire _06622_;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire net1738;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire net120;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire net1684;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire net1751;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire _06871_;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire _06875_;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire net1735;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire _06888_;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire net63;
 wire _06905_;
 wire _06906_;
 wire _06907_;
 wire net116;
 wire net115;
 wire _06910_;
 wire _06911_;
 wire net114;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire net113;
 wire _06922_;
 wire _06923_;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire _06939_;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire net62;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_26_clk;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire net1728;
 wire _06971_;
 wire net92;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire clknet_leaf_25_clk;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire net106;
 wire net105;
 wire net104;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire net103;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_0_clk;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire net141;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire net108;
 wire net107;
 wire net1916;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire net1918;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire net61;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire net60;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire \acc[0] ;
 wire \acc[10] ;
 wire \acc[11] ;
 wire \acc[12] ;
 wire \acc[13] ;
 wire \acc[14] ;
 wire \acc[15] ;
 wire \acc[1] ;
 wire \acc[2] ;
 wire \acc[3] ;
 wire \acc[4] ;
 wire \acc[5] ;
 wire \acc[6] ;
 wire \acc[7] ;
 wire \acc[8] ;
 wire \acc[9] ;
 wire \acc_sub.add_renorm0.exp[0] ;
 wire \acc_sub.add_renorm0.exp[1] ;
 wire \acc_sub.add_renorm0.exp[2] ;
 wire \acc_sub.add_renorm0.exp[3] ;
 wire \acc_sub.add_renorm0.exp[4] ;
 wire \acc_sub.add_renorm0.exp[5] ;
 wire \acc_sub.add_renorm0.exp[6] ;
 wire \acc_sub.add_renorm0.exp[7] ;
 wire \acc_sub.add_renorm0.mantisa[0] ;
 wire \acc_sub.add_renorm0.mantisa[10] ;
 wire \acc_sub.add_renorm0.mantisa[11] ;
 wire \acc_sub.add_renorm0.mantisa[1] ;
 wire \acc_sub.add_renorm0.mantisa[2] ;
 wire \acc_sub.add_renorm0.mantisa[3] ;
 wire \acc_sub.add_renorm0.mantisa[4] ;
 wire \acc_sub.add_renorm0.mantisa[5] ;
 wire \acc_sub.add_renorm0.mantisa[6] ;
 wire \acc_sub.add_renorm0.mantisa[7] ;
 wire \acc_sub.add_renorm0.mantisa[8] ;
 wire \acc_sub.add_renorm0.mantisa[9] ;
 wire \acc_sub.exp_mant_logic0.a[0] ;
 wire \acc_sub.exp_mant_logic0.a[10] ;
 wire \acc_sub.exp_mant_logic0.a[11] ;
 wire \acc_sub.exp_mant_logic0.a[12] ;
 wire \acc_sub.exp_mant_logic0.a[13] ;
 wire \acc_sub.exp_mant_logic0.a[14] ;
 wire \acc_sub.exp_mant_logic0.a[15] ;
 wire \acc_sub.exp_mant_logic0.a[1] ;
 wire \acc_sub.exp_mant_logic0.a[2] ;
 wire \acc_sub.exp_mant_logic0.a[3] ;
 wire \acc_sub.exp_mant_logic0.a[4] ;
 wire \acc_sub.exp_mant_logic0.a[5] ;
 wire \acc_sub.exp_mant_logic0.a[6] ;
 wire \acc_sub.exp_mant_logic0.a[7] ;
 wire \acc_sub.exp_mant_logic0.a[8] ;
 wire \acc_sub.exp_mant_logic0.a[9] ;
 wire \acc_sub.exp_mant_logic0.b[0] ;
 wire \acc_sub.exp_mant_logic0.b[10] ;
 wire \acc_sub.exp_mant_logic0.b[11] ;
 wire \acc_sub.exp_mant_logic0.b[12] ;
 wire \acc_sub.exp_mant_logic0.b[13] ;
 wire \acc_sub.exp_mant_logic0.b[14] ;
 wire \acc_sub.exp_mant_logic0.b[15] ;
 wire \acc_sub.exp_mant_logic0.b[1] ;
 wire \acc_sub.exp_mant_logic0.b[2] ;
 wire \acc_sub.exp_mant_logic0.b[3] ;
 wire \acc_sub.exp_mant_logic0.b[4] ;
 wire \acc_sub.exp_mant_logic0.b[5] ;
 wire \acc_sub.exp_mant_logic0.b[6] ;
 wire \acc_sub.exp_mant_logic0.b[7] ;
 wire \acc_sub.exp_mant_logic0.b[8] ;
 wire \acc_sub.exp_mant_logic0.b[9] ;
 wire \acc_sub.op_sign_logic0.add_sub ;
 wire \acc_sub.op_sign_logic0.mantisa_a[0] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[10] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[1] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[2] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[3] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[4] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[5] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[6] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[7] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[8] ;
 wire \acc_sub.op_sign_logic0.mantisa_a[9] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[0] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[10] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[1] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[2] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[3] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[4] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[5] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[6] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[7] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[8] ;
 wire \acc_sub.op_sign_logic0.mantisa_b[9] ;
 wire \acc_sub.op_sign_logic0.s_a ;
 wire \acc_sub.op_sign_logic0.s_b ;
 wire \acc_sub.reg1en.d[0] ;
 wire \acc_sub.reg1en.q[0] ;
 wire \acc_sub.reg2en.q[0] ;
 wire \acc_sub.reg3en.q[0] ;
 wire \acc_sub.reg4en.q[0] ;
 wire \acc_sub.reg_add_sub.q[0] ;
 wire \acc_sub.seg_reg0.q[22] ;
 wire \acc_sub.seg_reg0.q[23] ;
 wire \acc_sub.seg_reg0.q[24] ;
 wire \acc_sub.seg_reg0.q[25] ;
 wire \acc_sub.seg_reg0.q[26] ;
 wire \acc_sub.seg_reg0.q[27] ;
 wire \acc_sub.seg_reg0.q[28] ;
 wire \acc_sub.seg_reg0.q[29] ;
 wire \acc_sub.seg_reg1.q[20] ;
 wire \acc_sub.seg_reg1.q[21] ;
 wire \acc_sub.x2[0] ;
 wire \acc_sub.x2[10] ;
 wire \acc_sub.x2[11] ;
 wire \acc_sub.x2[12] ;
 wire \acc_sub.x2[13] ;
 wire \acc_sub.x2[14] ;
 wire \acc_sub.x2[15] ;
 wire \acc_sub.x2[1] ;
 wire \acc_sub.x2[2] ;
 wire \acc_sub.x2[3] ;
 wire \acc_sub.x2[4] ;
 wire \acc_sub.x2[5] ;
 wire \acc_sub.x2[6] ;
 wire \acc_sub.x2[7] ;
 wire \acc_sub.x2[8] ;
 wire \acc_sub.x2[9] ;
 wire \acc_sub.y[0] ;
 wire \acc_sub.y[10] ;
 wire \acc_sub.y[11] ;
 wire \acc_sub.y[12] ;
 wire \acc_sub.y[13] ;
 wire \acc_sub.y[14] ;
 wire \acc_sub.y[15] ;
 wire \acc_sub.y[1] ;
 wire \acc_sub.y[2] ;
 wire \acc_sub.y[3] ;
 wire \acc_sub.y[4] ;
 wire \acc_sub.y[5] ;
 wire \acc_sub.y[6] ;
 wire \acc_sub.y[7] ;
 wire \acc_sub.y[8] ;
 wire \acc_sub.y[9] ;
 wire \acc_sum.add_renorm0.exp[0] ;
 wire \acc_sum.add_renorm0.exp[1] ;
 wire \acc_sum.add_renorm0.exp[2] ;
 wire \acc_sum.add_renorm0.exp[3] ;
 wire \acc_sum.add_renorm0.exp[4] ;
 wire \acc_sum.add_renorm0.exp[5] ;
 wire \acc_sum.add_renorm0.exp[6] ;
 wire \acc_sum.add_renorm0.exp[7] ;
 wire \acc_sum.add_renorm0.mantisa[0] ;
 wire \acc_sum.add_renorm0.mantisa[10] ;
 wire \acc_sum.add_renorm0.mantisa[11] ;
 wire \acc_sum.add_renorm0.mantisa[1] ;
 wire \acc_sum.add_renorm0.mantisa[2] ;
 wire \acc_sum.add_renorm0.mantisa[3] ;
 wire \acc_sum.add_renorm0.mantisa[4] ;
 wire \acc_sum.add_renorm0.mantisa[5] ;
 wire \acc_sum.add_renorm0.mantisa[6] ;
 wire \acc_sum.add_renorm0.mantisa[7] ;
 wire \acc_sum.add_renorm0.mantisa[8] ;
 wire \acc_sum.add_renorm0.mantisa[9] ;
 wire \acc_sum.exp_mant_logic0.a[0] ;
 wire \acc_sum.exp_mant_logic0.a[10] ;
 wire \acc_sum.exp_mant_logic0.a[11] ;
 wire \acc_sum.exp_mant_logic0.a[12] ;
 wire \acc_sum.exp_mant_logic0.a[13] ;
 wire \acc_sum.exp_mant_logic0.a[14] ;
 wire \acc_sum.exp_mant_logic0.a[15] ;
 wire \acc_sum.exp_mant_logic0.a[1] ;
 wire \acc_sum.exp_mant_logic0.a[2] ;
 wire \acc_sum.exp_mant_logic0.a[3] ;
 wire \acc_sum.exp_mant_logic0.a[4] ;
 wire \acc_sum.exp_mant_logic0.a[5] ;
 wire \acc_sum.exp_mant_logic0.a[6] ;
 wire \acc_sum.exp_mant_logic0.a[7] ;
 wire \acc_sum.exp_mant_logic0.a[8] ;
 wire \acc_sum.exp_mant_logic0.a[9] ;
 wire \acc_sum.exp_mant_logic0.b[0] ;
 wire \acc_sum.exp_mant_logic0.b[10] ;
 wire \acc_sum.exp_mant_logic0.b[11] ;
 wire \acc_sum.exp_mant_logic0.b[12] ;
 wire \acc_sum.exp_mant_logic0.b[13] ;
 wire \acc_sum.exp_mant_logic0.b[14] ;
 wire \acc_sum.exp_mant_logic0.b[15] ;
 wire \acc_sum.exp_mant_logic0.b[1] ;
 wire \acc_sum.exp_mant_logic0.b[2] ;
 wire \acc_sum.exp_mant_logic0.b[3] ;
 wire \acc_sum.exp_mant_logic0.b[4] ;
 wire \acc_sum.exp_mant_logic0.b[5] ;
 wire \acc_sum.exp_mant_logic0.b[6] ;
 wire \acc_sum.exp_mant_logic0.b[7] ;
 wire \acc_sum.exp_mant_logic0.b[8] ;
 wire \acc_sum.exp_mant_logic0.b[9] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[0] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[10] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[1] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[2] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[3] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[4] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[5] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[6] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[7] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[8] ;
 wire \acc_sum.op_sign_logic0.mantisa_a[9] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[0] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[10] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[1] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[2] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[3] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[4] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[5] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[6] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[7] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[8] ;
 wire \acc_sum.op_sign_logic0.mantisa_b[9] ;
 wire \acc_sum.op_sign_logic0.s_a ;
 wire \acc_sum.op_sign_logic0.s_b ;
 wire \acc_sum.reg1en.d[0] ;
 wire \acc_sum.reg1en.q[0] ;
 wire \acc_sum.reg2en.q[0] ;
 wire \acc_sum.reg3en.q[0] ;
 wire \acc_sum.reg4en.q[0] ;
 wire \acc_sum.seg_reg0.q[22] ;
 wire \acc_sum.seg_reg0.q[23] ;
 wire \acc_sum.seg_reg0.q[24] ;
 wire \acc_sum.seg_reg0.q[25] ;
 wire \acc_sum.seg_reg0.q[26] ;
 wire \acc_sum.seg_reg0.q[27] ;
 wire \acc_sum.seg_reg0.q[28] ;
 wire \acc_sum.seg_reg0.q[29] ;
 wire \acc_sum.seg_reg1.q[20] ;
 wire \acc_sum.seg_reg1.q[21] ;
 wire \acc_sum.y[0] ;
 wire \acc_sum.y[10] ;
 wire \acc_sum.y[11] ;
 wire \acc_sum.y[12] ;
 wire \acc_sum.y[13] ;
 wire \acc_sum.y[14] ;
 wire \acc_sum.y[15] ;
 wire \acc_sum.y[1] ;
 wire \acc_sum.y[2] ;
 wire \acc_sum.y[3] ;
 wire \acc_sum.y[4] ;
 wire \acc_sum.y[5] ;
 wire \acc_sum.y[6] ;
 wire \acc_sum.y[7] ;
 wire \acc_sum.y[8] ;
 wire \acc_sum.y[9] ;
 wire \add_result[0] ;
 wire \add_result[10] ;
 wire \add_result[11] ;
 wire \add_result[12] ;
 wire \add_result[13] ;
 wire \add_result[14] ;
 wire \add_result[15] ;
 wire \add_result[1] ;
 wire \add_result[2] ;
 wire \add_result[3] ;
 wire \add_result[4] ;
 wire \add_result[5] ;
 wire \add_result[6] ;
 wire \add_result[7] ;
 wire \add_result[8] ;
 wire \add_result[9] ;
 wire \div_result[0] ;
 wire \div_result[10] ;
 wire \div_result[11] ;
 wire \div_result[12] ;
 wire \div_result[13] ;
 wire \div_result[14] ;
 wire \div_result[15] ;
 wire \div_result[1] ;
 wire \div_result[2] ;
 wire \div_result[3] ;
 wire \div_result[4] ;
 wire \div_result[5] ;
 wire \div_result[6] ;
 wire \div_result[7] ;
 wire \div_result[8] ;
 wire \div_result[9] ;
 wire \fp16_res_pipe.add_renorm0.exp[0] ;
 wire \fp16_res_pipe.add_renorm0.exp[1] ;
 wire \fp16_res_pipe.add_renorm0.exp[2] ;
 wire \fp16_res_pipe.add_renorm0.exp[3] ;
 wire \fp16_res_pipe.add_renorm0.exp[4] ;
 wire \fp16_res_pipe.add_renorm0.exp[5] ;
 wire \fp16_res_pipe.add_renorm0.exp[6] ;
 wire \fp16_res_pipe.add_renorm0.exp[7] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[0] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[10] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[11] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[1] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[2] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[3] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[4] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[5] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[6] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[7] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[8] ;
 wire \fp16_res_pipe.add_renorm0.mantisa[9] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[0] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[10] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[11] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[12] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[13] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[14] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[15] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[1] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[2] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[3] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[4] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[5] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[6] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[7] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[8] ;
 wire \fp16_res_pipe.exp_mant_logic0.a[9] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[0] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[10] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[11] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[12] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[13] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[14] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[15] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[1] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[2] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[3] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[4] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[5] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[6] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[7] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[8] ;
 wire \fp16_res_pipe.exp_mant_logic0.b[9] ;
 wire \fp16_res_pipe.op_sign_logic0.add_sub ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[0] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[10] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[1] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[2] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[3] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[4] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[5] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[6] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[7] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[8] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_a[9] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[0] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[10] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[1] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[2] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[3] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[4] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[5] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[6] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[7] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[8] ;
 wire \fp16_res_pipe.op_sign_logic0.mantisa_b[9] ;
 wire \fp16_res_pipe.op_sign_logic0.s_a ;
 wire \fp16_res_pipe.op_sign_logic0.s_b ;
 wire \fp16_res_pipe.reg1en.d[0] ;
 wire \fp16_res_pipe.reg1en.q[0] ;
 wire \fp16_res_pipe.reg2en.q[0] ;
 wire \fp16_res_pipe.reg3en.q[0] ;
 wire \fp16_res_pipe.reg4en.q[0] ;
 wire \fp16_res_pipe.reg_add_sub.q[0] ;
 wire \fp16_res_pipe.seg_reg0.q[22] ;
 wire \fp16_res_pipe.seg_reg0.q[23] ;
 wire \fp16_res_pipe.seg_reg0.q[24] ;
 wire \fp16_res_pipe.seg_reg0.q[25] ;
 wire \fp16_res_pipe.seg_reg0.q[26] ;
 wire \fp16_res_pipe.seg_reg0.q[27] ;
 wire \fp16_res_pipe.seg_reg0.q[28] ;
 wire \fp16_res_pipe.seg_reg0.q[29] ;
 wire \fp16_res_pipe.seg_reg1.q[20] ;
 wire \fp16_res_pipe.seg_reg1.q[21] ;
 wire \fp16_res_pipe.x2[0] ;
 wire \fp16_res_pipe.x2[10] ;
 wire \fp16_res_pipe.x2[11] ;
 wire \fp16_res_pipe.x2[12] ;
 wire \fp16_res_pipe.x2[13] ;
 wire \fp16_res_pipe.x2[14] ;
 wire \fp16_res_pipe.x2[15] ;
 wire \fp16_res_pipe.x2[1] ;
 wire \fp16_res_pipe.x2[2] ;
 wire \fp16_res_pipe.x2[3] ;
 wire \fp16_res_pipe.x2[4] ;
 wire \fp16_res_pipe.x2[5] ;
 wire \fp16_res_pipe.x2[6] ;
 wire \fp16_res_pipe.x2[7] ;
 wire \fp16_res_pipe.x2[8] ;
 wire \fp16_res_pipe.x2[9] ;
 wire \fp16_res_pipe.y[0] ;
 wire \fp16_res_pipe.y[10] ;
 wire \fp16_res_pipe.y[11] ;
 wire \fp16_res_pipe.y[12] ;
 wire \fp16_res_pipe.y[13] ;
 wire \fp16_res_pipe.y[14] ;
 wire \fp16_res_pipe.y[15] ;
 wire \fp16_res_pipe.y[1] ;
 wire \fp16_res_pipe.y[2] ;
 wire \fp16_res_pipe.y[3] ;
 wire \fp16_res_pipe.y[4] ;
 wire \fp16_res_pipe.y[5] ;
 wire \fp16_res_pipe.y[6] ;
 wire \fp16_res_pipe.y[7] ;
 wire \fp16_res_pipe.y[8] ;
 wire \fp16_res_pipe.y[9] ;
 wire \fp16_sum_pipe.add_renorm0.exp[0] ;
 wire \fp16_sum_pipe.add_renorm0.exp[1] ;
 wire \fp16_sum_pipe.add_renorm0.exp[2] ;
 wire \fp16_sum_pipe.add_renorm0.exp[3] ;
 wire \fp16_sum_pipe.add_renorm0.exp[4] ;
 wire \fp16_sum_pipe.add_renorm0.exp[5] ;
 wire \fp16_sum_pipe.add_renorm0.exp[6] ;
 wire \fp16_sum_pipe.add_renorm0.exp[7] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[0] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[10] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[11] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[1] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[2] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[3] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[4] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[5] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[6] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[7] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[8] ;
 wire \fp16_sum_pipe.add_renorm0.mantisa[9] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[0] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[10] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[11] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[12] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[13] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[14] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[15] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[1] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[2] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[3] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[4] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[5] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[6] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[7] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[8] ;
 wire \fp16_sum_pipe.exp_mant_logic0.a[9] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[0] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[10] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[11] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[12] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[13] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[14] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[15] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[1] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[2] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[3] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[4] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[5] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[6] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[7] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[8] ;
 wire \fp16_sum_pipe.exp_mant_logic0.b[9] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[0] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[10] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[1] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[2] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[3] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[4] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[5] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[6] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[7] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[8] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_a[9] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[0] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[10] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[1] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[2] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[3] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[4] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[5] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[6] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[7] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[8] ;
 wire \fp16_sum_pipe.op_sign_logic0.mantisa_b[9] ;
 wire \fp16_sum_pipe.op_sign_logic0.s_a ;
 wire \fp16_sum_pipe.op_sign_logic0.s_b ;
 wire \fp16_sum_pipe.reg1en.d[0] ;
 wire \fp16_sum_pipe.reg1en.q[0] ;
 wire \fp16_sum_pipe.reg2en.q[0] ;
 wire \fp16_sum_pipe.reg3en.q[0] ;
 wire \fp16_sum_pipe.reg4en.q[0] ;
 wire \fp16_sum_pipe.seg_reg0.q[22] ;
 wire \fp16_sum_pipe.seg_reg0.q[23] ;
 wire \fp16_sum_pipe.seg_reg0.q[24] ;
 wire \fp16_sum_pipe.seg_reg0.q[25] ;
 wire \fp16_sum_pipe.seg_reg0.q[26] ;
 wire \fp16_sum_pipe.seg_reg0.q[27] ;
 wire \fp16_sum_pipe.seg_reg0.q[28] ;
 wire \fp16_sum_pipe.seg_reg0.q[29] ;
 wire \fp16_sum_pipe.seg_reg1.q[20] ;
 wire \fp16_sum_pipe.seg_reg1.q[21] ;
 wire \fpdiv.div_out[0] ;
 wire \fpdiv.div_out[10] ;
 wire \fpdiv.div_out[11] ;
 wire \fpdiv.div_out[1] ;
 wire \fpdiv.div_out[2] ;
 wire \fpdiv.div_out[3] ;
 wire \fpdiv.div_out[4] ;
 wire \fpdiv.div_out[5] ;
 wire \fpdiv.div_out[6] ;
 wire \fpdiv.div_out[7] ;
 wire \fpdiv.div_out[8] ;
 wire \fpdiv.div_out[9] ;
 wire \fpdiv.divider0.counter[0] ;
 wire \fpdiv.divider0.counter[1] ;
 wire \fpdiv.divider0.counter[2] ;
 wire \fpdiv.divider0.counter[3] ;
 wire \fpdiv.divider0.dividend[10] ;
 wire \fpdiv.divider0.dividend[4] ;
 wire \fpdiv.divider0.dividend[5] ;
 wire \fpdiv.divider0.dividend[6] ;
 wire \fpdiv.divider0.dividend[7] ;
 wire \fpdiv.divider0.dividend[8] ;
 wire \fpdiv.divider0.dividend[9] ;
 wire \fpdiv.divider0.divisor[10] ;
 wire \fpdiv.divider0.divisor[4] ;
 wire \fpdiv.divider0.divisor[5] ;
 wire \fpdiv.divider0.divisor[6] ;
 wire \fpdiv.divider0.divisor[7] ;
 wire \fpdiv.divider0.divisor[8] ;
 wire \fpdiv.divider0.divisor[9] ;
 wire \fpdiv.divider0.divisor_reg[10] ;
 wire \fpdiv.divider0.divisor_reg[11] ;
 wire \fpdiv.divider0.divisor_reg[4] ;
 wire \fpdiv.divider0.divisor_reg[5] ;
 wire \fpdiv.divider0.divisor_reg[6] ;
 wire \fpdiv.divider0.divisor_reg[7] ;
 wire \fpdiv.divider0.divisor_reg[8] ;
 wire \fpdiv.divider0.divisor_reg[9] ;
 wire \fpdiv.divider0.en_r ;
 wire \fpdiv.divider0.remainder_reg[10] ;
 wire \fpdiv.divider0.remainder_reg[11] ;
 wire \fpdiv.divider0.remainder_reg[12] ;
 wire \fpdiv.divider0.remainder_reg[4] ;
 wire \fpdiv.divider0.remainder_reg[5] ;
 wire \fpdiv.divider0.remainder_reg[6] ;
 wire \fpdiv.divider0.remainder_reg[7] ;
 wire \fpdiv.divider0.remainder_reg[8] ;
 wire \fpdiv.divider0.remainder_reg[9] ;
 wire \fpdiv.divider0.state ;
 wire \fpdiv.reg1en.d[0] ;
 wire \fpdiv.reg1en.q[0] ;
 wire net77;
 wire \fpdiv.reg2en.q[0] ;
 wire \fpdiv.reg_a_out[10] ;
 wire \fpdiv.reg_a_out[11] ;
 wire \fpdiv.reg_a_out[12] ;
 wire \fpdiv.reg_a_out[13] ;
 wire \fpdiv.reg_a_out[14] ;
 wire \fpdiv.reg_a_out[15] ;
 wire \fpdiv.reg_a_out[7] ;
 wire \fpdiv.reg_a_out[8] ;
 wire \fpdiv.reg_a_out[9] ;
 wire \fpdiv.reg_b_out[10] ;
 wire \fpdiv.reg_b_out[11] ;
 wire \fpdiv.reg_b_out[12] ;
 wire \fpdiv.reg_b_out[13] ;
 wire \fpdiv.reg_b_out[14] ;
 wire \fpdiv.reg_b_out[15] ;
 wire \fpdiv.reg_b_out[7] ;
 wire \fpdiv.reg_b_out[8] ;
 wire \fpdiv.reg_b_out[9] ;
 wire \fpmul.reg1en.d[0] ;
 wire \fpmul.reg1en.q[0] ;
 wire \fpmul.reg2en.q[0] ;
 wire \fpmul.reg3en.q[0] ;
 wire \fpmul.reg_a_out[0] ;
 wire \fpmul.reg_a_out[10] ;
 wire \fpmul.reg_a_out[11] ;
 wire \fpmul.reg_a_out[12] ;
 wire \fpmul.reg_a_out[13] ;
 wire \fpmul.reg_a_out[14] ;
 wire \fpmul.reg_a_out[15] ;
 wire \fpmul.reg_a_out[1] ;
 wire \fpmul.reg_a_out[2] ;
 wire \fpmul.reg_a_out[3] ;
 wire \fpmul.reg_a_out[4] ;
 wire \fpmul.reg_a_out[5] ;
 wire \fpmul.reg_a_out[6] ;
 wire \fpmul.reg_a_out[7] ;
 wire \fpmul.reg_a_out[8] ;
 wire \fpmul.reg_a_out[9] ;
 wire \fpmul.reg_b_out[0] ;
 wire \fpmul.reg_b_out[10] ;
 wire \fpmul.reg_b_out[11] ;
 wire \fpmul.reg_b_out[12] ;
 wire \fpmul.reg_b_out[13] ;
 wire \fpmul.reg_b_out[14] ;
 wire \fpmul.reg_b_out[15] ;
 wire \fpmul.reg_b_out[1] ;
 wire \fpmul.reg_b_out[2] ;
 wire \fpmul.reg_b_out[3] ;
 wire \fpmul.reg_b_out[4] ;
 wire \fpmul.reg_b_out[5] ;
 wire \fpmul.reg_b_out[6] ;
 wire \fpmul.reg_b_out[7] ;
 wire \fpmul.reg_b_out[8] ;
 wire \fpmul.reg_b_out[9] ;
 wire \fpmul.reg_p_out[0] ;
 wire \fpmul.reg_p_out[10] ;
 wire \fpmul.reg_p_out[11] ;
 wire \fpmul.reg_p_out[12] ;
 wire \fpmul.reg_p_out[13] ;
 wire \fpmul.reg_p_out[14] ;
 wire \fpmul.reg_p_out[15] ;
 wire \fpmul.reg_p_out[1] ;
 wire \fpmul.reg_p_out[2] ;
 wire \fpmul.reg_p_out[3] ;
 wire \fpmul.reg_p_out[4] ;
 wire \fpmul.reg_p_out[5] ;
 wire \fpmul.reg_p_out[6] ;
 wire \fpmul.reg_p_out[7] ;
 wire \fpmul.reg_p_out[8] ;
 wire \fpmul.reg_p_out[9] ;
 wire \fpmul.result[15] ;
 wire \fpmul.seg_reg0.q[10] ;
 wire \fpmul.seg_reg0.q[11] ;
 wire \fpmul.seg_reg0.q[12] ;
 wire \fpmul.seg_reg0.q[13] ;
 wire \fpmul.seg_reg0.q[14] ;
 wire \fpmul.seg_reg0.q[15] ;
 wire \fpmul.seg_reg0.q[16] ;
 wire \fpmul.seg_reg0.q[17] ;
 wire \fpmul.seg_reg0.q[18] ;
 wire \fpmul.seg_reg0.q[19] ;
 wire \fpmul.seg_reg0.q[20] ;
 wire \fpmul.seg_reg0.q[21] ;
 wire \fpmul.seg_reg0.q[22] ;
 wire \fpmul.seg_reg0.q[23] ;
 wire \fpmul.seg_reg0.q[24] ;
 wire \fpmul.seg_reg0.q[25] ;
 wire \fpmul.seg_reg0.q[26] ;
 wire \fpmul.seg_reg0.q[27] ;
 wire \fpmul.seg_reg0.q[28] ;
 wire \fpmul.seg_reg0.q[29] ;
 wire \fpmul.seg_reg0.q[30] ;
 wire \fpmul.seg_reg0.q[31] ;
 wire \fpmul.seg_reg0.q[32] ;
 wire \fpmul.seg_reg0.q[33] ;
 wire \fpmul.seg_reg0.q[34] ;
 wire \fpmul.seg_reg0.q[35] ;
 wire \fpmul.seg_reg0.q[36] ;
 wire \fpmul.seg_reg0.q[37] ;
 wire \fpmul.seg_reg0.q[38] ;
 wire \fpmul.seg_reg0.q[39] ;
 wire \fpmul.seg_reg0.q[40] ;
 wire \fpmul.seg_reg0.q[41] ;
 wire \fpmul.seg_reg0.q[42] ;
 wire \fpmul.seg_reg0.q[43] ;
 wire \fpmul.seg_reg0.q[44] ;
 wire \fpmul.seg_reg0.q[45] ;
 wire \fpmul.seg_reg0.q[46] ;
 wire \fpmul.seg_reg0.q[47] ;
 wire \fpmul.seg_reg0.q[48] ;
 wire \fpmul.seg_reg0.q[49] ;
 wire \fpmul.seg_reg0.q[4] ;
 wire \fpmul.seg_reg0.q[50] ;
 wire \fpmul.seg_reg0.q[51] ;
 wire \fpmul.seg_reg0.q[52] ;
 wire \fpmul.seg_reg0.q[53] ;
 wire \fpmul.seg_reg0.q[5] ;
 wire \fpmul.seg_reg0.q[6] ;
 wire \fpmul.seg_reg0.q[7] ;
 wire \fpmul.seg_reg0.q[8] ;
 wire \fpmul.seg_reg0.q[9] ;
 wire \instr[0] ;
 wire \instr[10] ;
 wire \instr[11] ;
 wire \instr[12] ;
 wire \instr[13] ;
 wire \instr[14] ;
 wire \instr[15] ;
 wire \instr[1] ;
 wire \instr[2] ;
 wire \instr[3] ;
 wire \instr[4] ;
 wire \instr[5] ;
 wire \instr[6] ;
 wire \instr[7] ;
 wire \instr[8] ;
 wire \instr[9] ;
 wire load_en;
 wire net4;
 wire \piso.tx_active ;
 wire \piso.tx_bit_counter[0] ;
 wire \piso.tx_bit_counter[1] ;
 wire \piso.tx_bit_counter[2] ;
 wire \piso.tx_bit_counter[3] ;
 wire \piso.tx_bit_counter[4] ;
 wire \sipo.bit_counter[0] ;
 wire \sipo.bit_counter[1] ;
 wire \sipo.bit_counter[2] ;
 wire \sipo.bit_counter[3] ;
 wire \sipo.bit_counter[4] ;
 wire \sipo.receiving ;
 wire \sipo.shift_reg[10] ;
 wire \sipo.shift_reg[11] ;
 wire \sipo.shift_reg[12] ;
 wire \sipo.shift_reg[13] ;
 wire \sipo.shift_reg[14] ;
 wire \sipo.shift_reg[15] ;
 wire \sipo.shift_reg[1] ;
 wire \sipo.shift_reg[2] ;
 wire \sipo.shift_reg[3] ;
 wire \sipo.shift_reg[4] ;
 wire \sipo.shift_reg[5] ;
 wire \sipo.shift_reg[6] ;
 wire \sipo.shift_reg[7] ;
 wire \sipo.shift_reg[8] ;
 wire \sipo.shift_reg[9] ;
 wire \sipo.word[0] ;
 wire \sipo.word[10] ;
 wire \sipo.word[11] ;
 wire \sipo.word[12] ;
 wire \sipo.word[13] ;
 wire \sipo.word[14] ;
 wire \sipo.word[15] ;
 wire \sipo.word[1] ;
 wire \sipo.word[2] ;
 wire \sipo.word[3] ;
 wire \sipo.word[4] ;
 wire \sipo.word[5] ;
 wire \sipo.word[6] ;
 wire \sipo.word[7] ;
 wire \sipo.word[8] ;
 wire \sipo.word[9] ;
 wire \sipo.word_ready ;
 wire \state[0] ;
 wire \state[1] ;
 wire \state[2] ;
 wire \state[3] ;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1651;
 wire net1652;
 wire net1654;
 wire clknet_leaf_81_clk;
 wire net1647;
 wire net1648;
 wire net1669;
 wire clknet_leaf_89_clk;
 wire net1650;
 wire net1655;
 wire net1660;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_73_clk;
 wire net1659;
 wire net1662;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_53_clk;
 wire net1678;
 wire net1676;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_48_clk;
 wire net1686;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_40_clk;
 wire net1690;
 wire net1673;
 wire net1819;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_23_clk;
 wire net1685;
 wire net1677;
 wire clknet_leaf_32_clk;
 wire net1688;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_27_clk;
 wire net1687;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_6_clk;
 wire net1721;
 wire net1700;
 wire net140;
 wire net139;
 wire net138;
 wire net131;
 wire net1714;
 wire net1718;
 wire net1705;
 wire net1706;
 wire net1693;
 wire net128;
 wire net122;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1730;
 wire net112;
 wire net111;
 wire net1727;
 wire net1717;
 wire net1723;
 wire net1726;
 wire net1732;
 wire net1733;
 wire net1757;
 wire net102;
 wire net101;
 wire net1734;
 wire net98;
 wire net1762;
 wire net1740;
 wire net1742;
 wire net87;
 wire net1747;
 wire net1748;
 wire net83;
 wire net80;
 wire net1746;
 wire net1768;
 wire net1780;
 wire net73;
 wire net1894;
 wire net1817;
 wire net1766;
 wire net1758;
 wire net66;
 wire net1782;
 wire net1794;
 wire net1765;
 wire net1795;
 wire net1804;
 wire net1771;
 wire net1784;
 wire net1785;
 wire net1798;
 wire net1770;
 wire net54;
 wire net53;
 wire net1773;
 wire net1791;
 wire net1781;
 wire net1783;
 wire net1787;
 wire net1807;
 wire net1789;
 wire net47;
 wire net1803;
 wire net1850;
 wire net1778;
 wire net1800;
 wire net1806;
 wire net1827;
 wire net1805;
 wire net1796;
 wire net41;
 wire net43;
 wire net42;
 wire net44;
 wire net1797;
 wire net40;
 wire net1801;
 wire net1802;
 wire net1907;
 wire net1849;
 wire net1815;
 wire net1808;
 wire net1848;
 wire net1809;
 wire net1862;
 wire net1810;
 wire net1823;
 wire net1847;
 wire net1840;
 wire net1841;
 wire net1811;
 wire net1833;
 wire net1846;
 wire net1812;
 wire net1875;
 wire net1813;
 wire net1814;
 wire net1826;
 wire net1834;
 wire net1828;
 wire net1829;
 wire net1835;
 wire net1853;
 wire net1830;
 wire net38;
 wire net36;
 wire net37;
 wire net39;
 wire net1836;
 wire net1873;
 wire net1901;
 wire net1845;
 wire net1839;
 wire net1831;
 wire net1893;
 wire net34;
 wire net1852;
 wire net33;
 wire net35;
 wire net1832;
 wire net1837;
 wire net1838;
 wire net1872;
 wire net1842;
 wire net1871;
 wire net1843;
 wire net1854;
 wire net1917;
 wire net1892;
 wire net1844;
 wire net1874;
 wire net1905;
 wire net1900;
 wire net1890;
 wire net1915;
 wire net1855;
 wire net1913;
 wire net1912;
 wire net1902;
 wire net1914;
 wire net1891;
 wire net1923;
 wire net1932;
 wire net6;
 wire net2;
 wire net1909;
 wire net1945;
 wire net1910;
 wire net1953;
 wire net1856;
 wire net1899;
 wire net1857;
 wire net1858;
 wire net16;
 wire net1931;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1863;
 wire net1864;
 wire net1866;
 wire net1865;
 wire net1950;
 wire net17;
 wire net1867;
 wire net1928;
 wire net1868;
 wire net1930;
 wire net1869;
 wire net1929;
 wire net1870;
 wire net1920;
 wire net1925;
 wire net1946;
 wire net1927;
 wire net1952;
 wire net1933;
 wire net1937;
 wire net1942;
 wire net1938;
 wire net1939;
 wire net1934;
 wire net1940;
 wire net31;
 wire net1944;
 wire net1941;
 wire net30;
 wire net26;
 wire net27;
 wire net29;
 wire net28;
 wire net32;
 wire net1943;
 wire net1951;
 wire net1959;
 wire net1956;
 wire net1949;
 wire net15;
 wire net1958;
 wire net1962;
 wire net1954;
 wire net1961;
 wire net25;
 wire net7;
 wire net10;
 wire net1957;
 wire net1960;
 wire net9;
 wire net1;
 wire net3;
 wire net11;
 wire net1667;
 wire net8;
 wire net14;
 wire net13;
 wire net12;
 wire net1679;
 wire net1955;
 wire net1656;
 wire net1666;
 wire net1921;
 wire net1879;
 wire net1634;
 wire net1882;
 wire net1884;
 wire net23;
 wire net1883;
 wire net1878;
 wire net1880;
 wire net1877;
 wire net1881;
 wire net24;
 wire net1702;
 wire net1922;
 wire net1697;
 wire net1668;
 wire net1825;
 wire net1822;
 wire net21;
 wire net1779;
 wire net20;
 wire net1675;
 wire net1799;
 wire net1635;
 wire net19;
 wire net1786;
 wire net1680;
 wire net1696;
 wire net18;
 wire net22;
 wire net1897;
 wire net1935;
 wire net1729;
 wire net1720;
 wire net1695;
 wire net1681;
 wire net1636;
 wire net1948;
 wire net1896;
 wire net1777;
 wire net1924;
 wire net1898;
 wire net1926;
 wire net1947;
 wire net1903;
 wire net1904;
 wire net1936;
 wire net1699;
 wire net1637;
 wire net1682;
 wire net1895;
 wire net1911;
 wire net1908;
 wire net1906;
 wire net5;
 wire net1820;
 wire net1889;
 wire net1887;
 wire net1888;
 wire net1886;
 wire net1885;
 wire net1919;
 wire net1638;
 wire clknet_leaf_103_clk;
 wire clknet_leaf_104_clk;
 wire clknet_leaf_105_clk;
 wire clknet_leaf_106_clk;
 wire clknet_leaf_107_clk;
 wire clknet_leaf_108_clk;
 wire clknet_leaf_109_clk;
 wire clknet_leaf_110_clk;
 wire clknet_leaf_111_clk;
 wire clknet_leaf_112_clk;
 wire clknet_leaf_114_clk;
 wire clknet_leaf_115_clk;
 wire clknet_leaf_116_clk;
 wire clknet_leaf_117_clk;
 wire clknet_leaf_118_clk;
 wire clknet_leaf_119_clk;
 wire clknet_leaf_120_clk;
 wire clknet_leaf_121_clk;
 wire clknet_leaf_122_clk;
 wire clknet_leaf_123_clk;
 wire clknet_leaf_124_clk;
 wire clknet_leaf_125_clk;
 wire clknet_leaf_126_clk;
 wire clknet_leaf_127_clk;
 wire clknet_leaf_128_clk;
 wire clknet_leaf_129_clk;
 wire clknet_leaf_130_clk;
 wire clknet_leaf_131_clk;
 wire clknet_leaf_132_clk;
 wire clknet_leaf_134_clk;
 wire clknet_leaf_135_clk;
 wire clknet_leaf_136_clk;
 wire clknet_leaf_137_clk;
 wire clknet_leaf_139_clk;
 wire clknet_leaf_140_clk;
 wire clknet_leaf_141_clk;
 wire clknet_leaf_142_clk;
 wire clknet_leaf_143_clk;
 wire clknet_leaf_144_clk;
 wire clknet_0_clk;
 wire clknet_4_0_0_clk;
 wire clknet_4_1_0_clk;
 wire clknet_4_2_0_clk;
 wire clknet_4_3_0_clk;
 wire clknet_4_4_0_clk;
 wire clknet_4_5_0_clk;
 wire clknet_4_6_0_clk;
 wire clknet_4_7_0_clk;
 wire clknet_4_8_0_clk;
 wire clknet_4_9_0_clk;
 wire clknet_4_10_0_clk;
 wire clknet_4_11_0_clk;
 wire clknet_4_12_0_clk;
 wire clknet_4_13_0_clk;
 wire clknet_4_14_0_clk;
 wire clknet_4_15_0_clk;
 wire clknet_5_0__leaf_clk;
 wire clknet_5_1__leaf_clk;
 wire clknet_5_2__leaf_clk;
 wire clknet_5_3__leaf_clk;
 wire clknet_5_4__leaf_clk;
 wire clknet_5_5__leaf_clk;
 wire clknet_5_6__leaf_clk;
 wire clknet_5_7__leaf_clk;
 wire clknet_5_8__leaf_clk;
 wire clknet_5_9__leaf_clk;
 wire clknet_5_10__leaf_clk;
 wire clknet_5_11__leaf_clk;
 wire clknet_5_12__leaf_clk;
 wire clknet_5_13__leaf_clk;
 wire clknet_5_14__leaf_clk;
 wire clknet_5_15__leaf_clk;
 wire clknet_5_16__leaf_clk;
 wire clknet_5_17__leaf_clk;
 wire clknet_5_18__leaf_clk;
 wire clknet_5_19__leaf_clk;
 wire clknet_5_20__leaf_clk;
 wire clknet_5_21__leaf_clk;
 wire clknet_5_22__leaf_clk;
 wire clknet_5_23__leaf_clk;
 wire clknet_5_24__leaf_clk;
 wire clknet_5_25__leaf_clk;
 wire clknet_5_26__leaf_clk;
 wire clknet_5_27__leaf_clk;
 wire clknet_5_28__leaf_clk;
 wire clknet_5_29__leaf_clk;
 wire clknet_5_30__leaf_clk;
 wire clknet_5_31__leaf_clk;

 sg13g2_inv_2 _07117_ (.Y(_01490_),
    .A(\acc_sub.seg_reg1.q[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1821 (.A(\fp16_res_pipe.seg_reg1.q[21] ),
    .X(net1821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07119_ (.VDD(VPWR),
    .Y(_01492_),
    .A(\acc_sub.reg2en.q[0] ),
    .VSS(VGND));
 sg13g2_buf_2 place1816 (.A(\acc_sum.reg2en.q[0] ),
    .X(net1816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07121_ (.Y(_01494_),
    .A(\acc_sub.op_sign_logic0.s_a ),
    .B(\acc_sub.op_sign_logic0.s_b ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07122_ (.Y(_01495_),
    .A(\acc_sub.op_sign_logic0.add_sub ),
    .B(_01494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07123_ (.A(net1783),
    .B(_01495_),
    .Y(_01496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout74 (.A(net76),
    .X(net74),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07125_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01490_),
    .A2(_01492_),
    .Y(_01489_),
    .B1(_01496_));
 sg13g2_inv_1 _07126_ (.VDD(VPWR),
    .Y(_01498_),
    .A(\acc_sub.seg_reg1.q[20] ),
    .VSS(VGND));
 sg13g2_inv_1 _07127_ (.VDD(VPWR),
    .Y(_01499_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07128_ (.A(\acc_sub.op_sign_logic0.mantisa_b[10] ),
    .B(_01499_),
    .Y(_01500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07129_ (.VDD(VPWR),
    .Y(_01501_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07130_ (.A(\acc_sub.op_sign_logic0.mantisa_a[10] ),
    .B(_01501_),
    .Y(_01502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07131_ (.VDD(VPWR),
    .Y(_01503_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[8] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07132_ (.A(\acc_sub.op_sign_logic0.mantisa_b[8] ),
    .B(_01503_),
    .Y(_01504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07133_ (.VDD(VPWR),
    .Y(_01505_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[8] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07134_ (.A(\acc_sub.op_sign_logic0.mantisa_a[8] ),
    .B(_01505_),
    .Y(_01506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07135_ (.A(_01504_),
    .B(_01506_),
    .Y(_01507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07136_ (.VDD(VPWR),
    .Y(_01508_),
    .A(_01507_),
    .VSS(VGND));
 sg13g2_inv_1 _07137_ (.VDD(VPWR),
    .Y(_01509_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[9] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07138_ (.A(\acc_sub.op_sign_logic0.mantisa_b[9] ),
    .B(_01509_),
    .Y(_01510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07139_ (.Y(_01511_),
    .A(_01509_),
    .B(\acc_sub.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07140_ (.VDD(VPWR),
    .Y(_01512_),
    .A(_01511_),
    .VSS(VGND));
 sg13g2_nor2_2 _07141_ (.A(_01510_),
    .B(_01512_),
    .Y(_01513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07142_ (.VDD(VPWR),
    .Y(_01514_),
    .A(_01513_),
    .VSS(VGND));
 sg13g2_nor2_1 _07143_ (.A(_01508_),
    .B(_01514_),
    .Y(_01515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07144_ (.VDD(VPWR),
    .Y(_01516_),
    .A(_01515_),
    .VSS(VGND));
 sg13g2_inv_1 _07145_ (.VDD(VPWR),
    .Y(_01517_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07146_ (.A(\acc_sub.op_sign_logic0.mantisa_b[7] ),
    .B(_01517_),
    .Y(_01518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07147_ (.VDD(VPWR),
    .Y(_01519_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07148_ (.A(\acc_sub.op_sign_logic0.mantisa_a[7] ),
    .B(_01519_),
    .Y(_01520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07149_ (.A(_01518_),
    .B(_01520_),
    .Y(_01521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07150_ (.VDD(VPWR),
    .Y(_01522_),
    .A(_01521_),
    .VSS(VGND));
 sg13g2_inv_1 _07151_ (.VDD(VPWR),
    .Y(_01523_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[6] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07152_ (.A(\acc_sub.op_sign_logic0.mantisa_b[6] ),
    .B(_01523_),
    .Y(_01524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07153_ (.VDD(VPWR),
    .Y(_01525_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[6] ),
    .VSS(VGND));
 sg13g2_nor2_2 _07154_ (.A(\acc_sub.op_sign_logic0.mantisa_a[6] ),
    .B(_01525_),
    .Y(_01526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07155_ (.A(_01524_),
    .B(_01526_),
    .Y(_01527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07156_ (.VDD(VPWR),
    .Y(_01528_),
    .A(_01527_),
    .VSS(VGND));
 sg13g2_nor2_1 _07157_ (.A(_01522_),
    .B(_01528_),
    .Y(_01529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07158_ (.VDD(VPWR),
    .Y(_01530_),
    .A(_01529_),
    .VSS(VGND));
 sg13g2_inv_1 _07159_ (.VDD(VPWR),
    .Y(_01531_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07160_ (.A(\acc_sub.op_sign_logic0.mantisa_b[5] ),
    .B(_01531_),
    .Y(_01532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07161_ (.VDD(VPWR),
    .Y(_01533_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07162_ (.A(\acc_sub.op_sign_logic0.mantisa_a[5] ),
    .B(_01533_),
    .Y(_01534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07163_ (.A(_01532_),
    .B(_01534_),
    .Y(_01535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07164_ (.VDD(VPWR),
    .Y(_01536_),
    .A(_01535_),
    .VSS(VGND));
 sg13g2_inv_1 _07165_ (.VDD(VPWR),
    .Y(_01537_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[4] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07166_ (.A(\acc_sub.op_sign_logic0.mantisa_b[4] ),
    .B(_01537_),
    .Y(_01538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07167_ (.VDD(VPWR),
    .Y(_01539_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[4] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07168_ (.A(\acc_sub.op_sign_logic0.mantisa_a[4] ),
    .B(_01539_),
    .Y(_01540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07169_ (.A(_01538_),
    .B(_01540_),
    .Y(_01541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07170_ (.VDD(VPWR),
    .Y(_01542_),
    .A(_01541_),
    .VSS(VGND));
 sg13g2_nor2_1 _07171_ (.A(_01536_),
    .B(_01542_),
    .Y(_01543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07172_ (.VDD(VPWR),
    .Y(_01544_),
    .A(_01543_),
    .VSS(VGND));
 sg13g2_inv_1 _07173_ (.VDD(VPWR),
    .Y(_01545_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[0] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07174_ (.A(\acc_sub.op_sign_logic0.mantisa_a[0] ),
    .B(_01545_),
    .Y(_01546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07175_ (.VDD(VPWR),
    .Y(_01547_),
    .A(_01546_),
    .VSS(VGND));
 sg13g2_inv_1 _07176_ (.VDD(VPWR),
    .Y(_01548_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07177_ (.Y(_01549_),
    .A(_01548_),
    .B(\acc_sub.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07178_ (.VDD(VPWR),
    .Y(_01550_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07179_ (.Y(_01551_),
    .A(_01550_),
    .B(\acc_sub.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07180_ (.VDD(VPWR),
    .Y(_01552_),
    .A(_01551_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01547_),
    .A2(_01549_),
    .Y(_01553_),
    .B1(_01552_));
 sg13g2_inv_1 _07182_ (.VDD(VPWR),
    .Y(_01554_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07183_ (.A(\acc_sub.op_sign_logic0.mantisa_a[3] ),
    .B(_01554_),
    .Y(_01555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07184_ (.VDD(VPWR),
    .Y(_01556_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07185_ (.A(\acc_sub.op_sign_logic0.mantisa_b[3] ),
    .B(_01556_),
    .Y(_01557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07186_ (.A(_01555_),
    .B(_01557_),
    .Y(_01558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07187_ (.Y(_01559_),
    .A(_01558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07188_ (.VDD(VPWR),
    .Y(_01560_),
    .A(\acc_sub.op_sign_logic0.mantisa_b[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07189_ (.A(\acc_sub.op_sign_logic0.mantisa_a[2] ),
    .B(_01560_),
    .Y(_01561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07190_ (.VDD(VPWR),
    .Y(_01562_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07191_ (.A(\acc_sub.op_sign_logic0.mantisa_b[2] ),
    .B(_01562_),
    .Y(_01563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07192_ (.A(_01561_),
    .B(_01563_),
    .Y(_01564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07193_ (.VDD(VPWR),
    .Y(_01565_),
    .A(_01564_),
    .VSS(VGND));
 sg13g2_nor2_1 _07194_ (.A(_01559_),
    .B(_01565_),
    .Y(_01566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07195_ (.VDD(VPWR),
    .Y(_01567_),
    .A(_01566_),
    .VSS(VGND));
 sg13g2_inv_1 _07196_ (.VDD(VPWR),
    .Y(_01568_),
    .A(_01555_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07197_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01568_),
    .A2(_01563_),
    .Y(_01569_),
    .B1(_01557_));
 sg13g2_o21ai_1 _07198_ (.B1(_01569_),
    .VDD(VPWR),
    .Y(_01570_),
    .VSS(VGND),
    .A1(_01553_),
    .A2(_01567_));
 sg13g2_inv_1 _07199_ (.VDD(VPWR),
    .Y(_01571_),
    .A(_01570_),
    .VSS(VGND));
 sg13g2_inv_1 _07200_ (.VDD(VPWR),
    .Y(_01572_),
    .A(_01534_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07201_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01572_),
    .A2(_01538_),
    .Y(_01573_),
    .B1(_01532_));
 sg13g2_o21ai_1 _07202_ (.B1(_01573_),
    .VDD(VPWR),
    .Y(_01574_),
    .VSS(VGND),
    .A1(_01544_),
    .A2(_01571_));
 sg13g2_inv_1 _07203_ (.VDD(VPWR),
    .Y(_01575_),
    .A(_01574_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07204_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01521_),
    .A2(_01524_),
    .Y(_01576_),
    .B1(_01518_));
 sg13g2_o21ai_1 _07205_ (.B1(_01576_),
    .VDD(VPWR),
    .Y(_01577_),
    .VSS(VGND),
    .A1(_01530_),
    .A2(_01575_));
 sg13g2_inv_1 _07206_ (.VDD(VPWR),
    .Y(_01578_),
    .A(_01577_),
    .VSS(VGND));
 sg13g2_o21ai_1 _07207_ (.B1(_01511_),
    .VDD(VPWR),
    .Y(_01579_),
    .VSS(VGND),
    .A1(_01510_),
    .A2(_01504_));
 sg13g2_o21ai_1 _07208_ (.B1(_01579_),
    .VDD(VPWR),
    .Y(_01580_),
    .VSS(VGND),
    .A1(_01516_),
    .A2(_01578_));
 sg13g2_nor2_1 _07209_ (.A(_01530_),
    .B(_01516_),
    .Y(_01581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07210_ (.Y(_01582_),
    .A(_01551_),
    .B(_01549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07211_ (.A(_01500_),
    .B(_01502_),
    .Y(_01583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07212_ (.VDD(VPWR),
    .Y(_01584_),
    .A(_01583_),
    .VSS(VGND));
 sg13g2_nor2b_1 _07213_ (.A(\acc_sub.op_sign_logic0.mantisa_b[0] ),
    .B_N(\acc_sub.op_sign_logic0.mantisa_a[0] ),
    .Y(_01585_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07214_ (.VDD(VPWR),
    .Y(_01586_),
    .A(_01585_),
    .VSS(VGND));
 sg13g2_nand2_1 _07215_ (.Y(_01587_),
    .A(_01586_),
    .B(_01547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07216_ (.A(_01582_),
    .B(_01584_),
    .C(_01587_),
    .Y(_01588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _07217_ (.B(_01543_),
    .C(_01566_),
    .A(_01581_),
    .Y(_01589_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01588_));
 sg13g2_nand3b_1 _07218_ (.B(_01580_),
    .C(_01589_),
    .Y(_01590_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_01502_));
 sg13g2_nor2b_2 _07219_ (.A(_01500_),
    .B_N(_01590_),
    .Y(_01591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_46_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_46_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07222_ (.Y(_01594_),
    .A(\acc_sub.op_sign_logic0.s_b ),
    .B(\acc_sub.op_sign_logic0.add_sub ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07223_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01591_),
    .A2(_01594_),
    .Y(_01595_),
    .B1(_01492_));
 sg13g2_o21ai_1 _07224_ (.B1(_01595_),
    .VDD(VPWR),
    .Y(_01596_),
    .VSS(VGND),
    .A1(\acc_sub.op_sign_logic0.s_a ),
    .A2(_01591_));
 sg13g2_o21ai_1 _07225_ (.B1(_01596_),
    .VDD(VPWR),
    .Y(_01488_),
    .VSS(VGND),
    .A1(net1798),
    .A2(_01498_));
 sg13g2_nand2_1 _07226_ (.Y(_01597_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[0] ),
    .B(\acc_sub.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07227_ (.Y(_01598_),
    .B(_01582_),
    .A_N(_01597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07228_ (.B1(_01598_),
    .VDD(VPWR),
    .Y(_01599_),
    .VSS(VGND),
    .A1(_01548_),
    .A2(_01550_));
 sg13g2_nand2_1 _07229_ (.Y(_01600_),
    .A(_01599_),
    .B(_01565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07230_ (.B1(_01600_),
    .VDD(VPWR),
    .Y(_01601_),
    .VSS(VGND),
    .A1(_01562_),
    .A2(_01560_));
 sg13g2_nand2_1 _07231_ (.Y(_01602_),
    .A(_01601_),
    .B(_01559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07232_ (.B1(_01602_),
    .VDD(VPWR),
    .Y(_01603_),
    .VSS(VGND),
    .A1(_01556_),
    .A2(_01554_));
 sg13g2_nand2_1 _07233_ (.Y(_01604_),
    .A(_01603_),
    .B(_01542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07234_ (.B1(_01604_),
    .VDD(VPWR),
    .Y(_01605_),
    .VSS(VGND),
    .A1(_01537_),
    .A2(_01539_));
 sg13g2_nand2_1 _07235_ (.Y(_01606_),
    .A(_01605_),
    .B(_01536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07236_ (.B1(_01606_),
    .VDD(VPWR),
    .Y(_01607_),
    .VSS(VGND),
    .A1(_01531_),
    .A2(_01533_));
 sg13g2_nand2_1 _07237_ (.Y(_01608_),
    .A(_01607_),
    .B(_01528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07238_ (.B1(_01608_),
    .VDD(VPWR),
    .Y(_01609_),
    .VSS(VGND),
    .A1(_01523_),
    .A2(_01525_));
 sg13g2_nand2_1 _07239_ (.Y(_01610_),
    .A(_01609_),
    .B(_01522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07240_ (.B1(_01610_),
    .VDD(VPWR),
    .Y(_01611_),
    .VSS(VGND),
    .A1(_01517_),
    .A2(_01519_));
 sg13g2_nand2_1 _07241_ (.Y(_01612_),
    .A(_01611_),
    .B(_01508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07242_ (.B1(_01612_),
    .VDD(VPWR),
    .Y(_01613_),
    .VSS(VGND),
    .A1(_01503_),
    .A2(_01505_));
 sg13g2_nand2_1 _07243_ (.Y(_01614_),
    .A(_01613_),
    .B(_01514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07244_ (.Y(_01615_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[9] ),
    .B(\acc_sub.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07245_ (.A2(_01615_),
    .A1(_01614_),
    .B1(_01583_),
    .X(_01616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07246_ (.B1(_01616_),
    .VDD(VPWR),
    .Y(_01617_),
    .VSS(VGND),
    .A1(_01499_),
    .A2(_01501_));
 sg13g2_nand2_1 _07247_ (.Y(_01618_),
    .A(_01617_),
    .B(_01496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07248_ (.Y(_01619_),
    .A(net1784),
    .B(\acc_sub.add_renorm0.mantisa[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07249_ (.Y(_01487_),
    .A(_01618_),
    .B(_01619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07250_ (.B(_01583_),
    .C(_01615_),
    .A(_01614_),
    .Y(_01620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07251_ (.B(_01620_),
    .C(net1744),
    .A(_01616_),
    .Y(_01621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07252_ (.Y(_01622_),
    .A(net1783),
    .B(\acc_sub.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07253_ (.VDD(VPWR),
    .Y(_01623_),
    .A(_01549_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07254_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01586_),
    .A2(_01551_),
    .Y(_01624_),
    .B1(_01623_));
 sg13g2_inv_1 _07255_ (.VDD(VPWR),
    .Y(_01625_),
    .A(_01624_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07256_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01625_),
    .A2(_01564_),
    .Y(_01626_),
    .B1(_01561_));
 sg13g2_a21oi_1 _07257_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01626_),
    .A2(_01568_),
    .Y(_01627_),
    .B1(_01557_));
 sg13g2_a21oi_1 _07258_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01627_),
    .A2(_01541_),
    .Y(_01628_),
    .B1(_01540_));
 sg13g2_a21oi_1 _07259_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01628_),
    .A2(_01572_),
    .Y(_01629_),
    .B1(_01532_));
 sg13g2_inv_1 _07260_ (.VDD(VPWR),
    .Y(_01630_),
    .A(_01629_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07261_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01521_),
    .A2(_01526_),
    .Y(_01631_),
    .B1(_01520_));
 sg13g2_o21ai_1 _07262_ (.B1(_01631_),
    .VDD(VPWR),
    .Y(_01632_),
    .VSS(VGND),
    .A1(_01530_),
    .A2(_01630_));
 sg13g2_a221oi_1 _07263_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01515_),
    .C1(_01512_),
    .B1(_01632_),
    .A1(_01506_),
    .Y(_01633_),
    .A2(_01513_));
 sg13g2_o21ai_1 _07264_ (.B1(_01590_),
    .VDD(VPWR),
    .Y(_01634_),
    .VSS(VGND),
    .A1(_01500_),
    .A2(_01633_));
 sg13g2_inv_1 _07265_ (.VDD(VPWR),
    .Y(_01635_),
    .A(_01495_),
    .VSS(VGND));
 sg13g2_nor2_2 _07266_ (.A(net1783),
    .B(_01635_),
    .Y(_01636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07267_ (.B(_01636_),
    .C(_01584_),
    .A(_01634_),
    .Y(_01637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07268_ (.B(_01622_),
    .C(_01637_),
    .A(_01621_),
    .Y(_01486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07269_ (.Y(_01638_),
    .B(_01513_),
    .A_N(_01613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07270_ (.B(net1744),
    .C(_01614_),
    .A(_01638_),
    .Y(_01639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07271_ (.Y(_01640_),
    .A(net1783),
    .B(\acc_sub.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _07272_ (.A2(_01507_),
    .A1(_01577_),
    .B1(_01504_),
    .X(_01641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01632_),
    .A2(_01507_),
    .Y(_01642_),
    .B1(_01506_));
 sg13g2_nand2_1 _07274_ (.Y(_01643_),
    .A(net1665),
    .B(_01642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07275_ (.B1(_01643_),
    .VDD(VPWR),
    .Y(_01644_),
    .VSS(VGND),
    .A1(net1665),
    .A2(_01641_));
 sg13g2_xnor2_1 _07276_ (.Y(_01645_),
    .A(_01513_),
    .B(_01644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07277_ (.Y(_01646_),
    .A(_01645_),
    .B(_01636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07278_ (.B(_01640_),
    .C(_01646_),
    .A(_01639_),
    .Y(_01485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07279_ (.Y(_01647_),
    .A(\acc_sub.add_renorm0.mantisa[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07280_ (.A(_01508_),
    .B(_01611_),
    .Y(_01648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07281_ (.VDD(VPWR),
    .Y(_01649_),
    .A(_01612_),
    .VSS(VGND));
 sg13g2_nor3_1 _07282_ (.A(net1783),
    .B(_01648_),
    .C(_01649_),
    .Y(_01650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07283_ (.A(_01578_),
    .B(net1665),
    .Y(_01651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07284_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01632_),
    .A2(net1665),
    .Y(_01652_),
    .B1(_01651_));
 sg13g2_a21oi_1 _07285_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01652_),
    .A2(_01507_),
    .Y(_01653_),
    .B1(_01635_));
 sg13g2_o21ai_1 _07286_ (.B1(_01653_),
    .VDD(VPWR),
    .Y(_01654_),
    .VSS(VGND),
    .A1(_01507_),
    .A2(_01652_));
 sg13g2_o21ai_1 _07287_ (.B1(_01654_),
    .VDD(VPWR),
    .Y(_01655_),
    .VSS(VGND),
    .A1(_01636_),
    .A2(_01650_));
 sg13g2_o21ai_1 _07288_ (.B1(_01655_),
    .VDD(VPWR),
    .Y(_01484_),
    .VSS(VGND),
    .A1(\acc_sub.reg2en.q[0] ),
    .A2(_01647_));
 sg13g2_inv_2 _07289_ (.Y(_01656_),
    .A(_01636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07290_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01574_),
    .A2(_01527_),
    .Y(_01657_),
    .B1(_01524_));
 sg13g2_nor2_1 _07291_ (.A(_01528_),
    .B(_01630_),
    .Y(_01658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07292_ (.B1(net1667),
    .VDD(VPWR),
    .Y(_01659_),
    .VSS(VGND),
    .A1(_01526_),
    .A2(_01658_));
 sg13g2_o21ai_1 _07293_ (.B1(_01659_),
    .VDD(VPWR),
    .Y(_01660_),
    .VSS(VGND),
    .A1(net1667),
    .A2(_01657_));
 sg13g2_xnor2_1 _07294_ (.Y(_01661_),
    .A(_01521_),
    .B(_01660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07295_ (.Y(_01662_),
    .A(_01521_),
    .B(_01609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07296_ (.Y(_01663_),
    .B1(net1744),
    .B2(_01662_),
    .A2(\acc_sub.add_renorm0.mantisa[7] ),
    .A1(net1784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07297_ (.B1(_01663_),
    .VDD(VPWR),
    .Y(_01483_),
    .VSS(VGND),
    .A1(_01656_),
    .A2(_01661_));
 sg13g2_nand2_1 _07298_ (.Y(_01664_),
    .A(net1667),
    .B(_01629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07299_ (.B1(_01664_),
    .VDD(VPWR),
    .Y(_01665_),
    .VSS(VGND),
    .A1(_01575_),
    .A2(net1667));
 sg13g2_a21oi_1 _07300_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01665_),
    .A2(_01527_),
    .Y(_01666_),
    .B1(_01656_));
 sg13g2_o21ai_1 _07301_ (.B1(_01666_),
    .VDD(VPWR),
    .Y(_01667_),
    .VSS(VGND),
    .A1(_01527_),
    .A2(_01665_));
 sg13g2_nand2_1 _07302_ (.Y(_01668_),
    .A(net1784),
    .B(\acc_sub.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07303_ (.Y(_01669_),
    .B(_01527_),
    .A_N(_01607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07304_ (.B(net1744),
    .C(_01608_),
    .A(_01669_),
    .Y(_01670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07305_ (.B(_01668_),
    .C(_01670_),
    .A(_01667_),
    .Y(_01482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07306_ (.A(_01542_),
    .B(_01571_),
    .Y(_01671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07307_ (.A(_01538_),
    .B(_01671_),
    .C(net1667),
    .Y(_01672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07308_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01628_),
    .A2(net1667),
    .Y(_01673_),
    .B1(_01672_));
 sg13g2_xnor2_1 _07309_ (.Y(_01674_),
    .A(_01535_),
    .B(_01673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07310_ (.Y(_01675_),
    .A(_01535_),
    .B(_01605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07311_ (.Y(_01676_),
    .B1(net1744),
    .B2(_01675_),
    .A2(\acc_sub.add_renorm0.mantisa[5] ),
    .A1(net1784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07312_ (.B1(_01676_),
    .VDD(VPWR),
    .Y(_01481_),
    .VSS(VGND),
    .A1(_01656_),
    .A2(_01674_));
 sg13g2_nand2_1 _07313_ (.Y(_01677_),
    .A(net1667),
    .B(_01627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07314_ (.B1(_01677_),
    .VDD(VPWR),
    .Y(_01678_),
    .VSS(VGND),
    .A1(_01571_),
    .A2(net1667));
 sg13g2_a21oi_1 _07315_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01678_),
    .A2(_01541_),
    .Y(_01679_),
    .B1(_01656_));
 sg13g2_o21ai_1 _07316_ (.B1(_01679_),
    .VDD(VPWR),
    .Y(_01680_),
    .VSS(VGND),
    .A1(_01541_),
    .A2(_01678_));
 sg13g2_nand2_1 _07317_ (.Y(_01681_),
    .A(net1784),
    .B(\acc_sub.add_renorm0.mantisa[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07318_ (.Y(_01682_),
    .B(_01541_),
    .A_N(_01603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07319_ (.B(net1744),
    .C(_01604_),
    .A(_01682_),
    .Y(_01683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07320_ (.B(_01681_),
    .C(_01683_),
    .A(_01680_),
    .Y(_01480_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07321_ (.VDD(VPWR),
    .Y(_01684_),
    .A(_01563_),
    .VSS(VGND));
 sg13g2_o21ai_1 _07322_ (.B1(_01684_),
    .VDD(VPWR),
    .Y(_01685_),
    .VSS(VGND),
    .A1(_01561_),
    .A2(_01553_));
 sg13g2_nand2_1 _07323_ (.Y(_01686_),
    .A(net1666),
    .B(_01626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07324_ (.B1(_01686_),
    .VDD(VPWR),
    .Y(_01687_),
    .VSS(VGND),
    .A1(net1666),
    .A2(_01685_));
 sg13g2_a21oi_1 _07325_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01687_),
    .A2(_01559_),
    .Y(_01688_),
    .B1(_01656_));
 sg13g2_o21ai_1 _07326_ (.B1(_01688_),
    .VDD(VPWR),
    .Y(_01689_),
    .VSS(VGND),
    .A1(_01559_),
    .A2(_01687_));
 sg13g2_nand2_1 _07327_ (.Y(_01690_),
    .A(net1784),
    .B(\acc_sub.add_renorm0.mantisa[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07328_ (.Y(_01691_),
    .B(_01558_),
    .A_N(_01601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07329_ (.B(net1744),
    .C(_01602_),
    .A(_01691_),
    .Y(_01692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07330_ (.B(_01690_),
    .C(_01692_),
    .A(_01689_),
    .Y(_01479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07331_ (.Y(_01693_),
    .A(net1666),
    .B(_01625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07332_ (.B1(_01693_),
    .VDD(VPWR),
    .Y(_01694_),
    .VSS(VGND),
    .A1(_01553_),
    .A2(net1666));
 sg13g2_and2_1 _07333_ (.A(_01694_),
    .B(_01564_),
    .X(_01695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07334_ (.B1(_01636_),
    .VDD(VPWR),
    .Y(_01696_),
    .VSS(VGND),
    .A1(_01564_),
    .A2(_01694_));
 sg13g2_nand2b_1 _07335_ (.Y(_01697_),
    .B(_01564_),
    .A_N(_01599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _07336_ (.A(_01600_),
    .B(net1744),
    .X(_01698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07337_ (.Y(_01699_),
    .B1(_01697_),
    .B2(_01698_),
    .A2(\acc_sub.add_renorm0.mantisa[2] ),
    .A1(net1784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07338_ (.B1(_01699_),
    .VDD(VPWR),
    .Y(_01478_),
    .VSS(VGND),
    .A1(_01695_),
    .A2(_01696_));
 sg13g2_inv_1 _07339_ (.VDD(VPWR),
    .Y(_01700_),
    .A(\acc_sub.add_renorm0.mantisa[1] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _07340_ (.Y(_01701_),
    .A(_01597_),
    .B(_01582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07341_ (.Y(_01702_),
    .A(net1665),
    .B(_01586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07342_ (.B1(_01702_),
    .VDD(VPWR),
    .Y(_01703_),
    .VSS(VGND),
    .A1(_01546_),
    .A2(net1665));
 sg13g2_xor2_1 _07343_ (.B(_01703_),
    .A(_01582_),
    .X(_01704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07344_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01704_),
    .A2(_01495_),
    .Y(_01705_),
    .B1(net1783));
 sg13g2_o21ai_1 _07345_ (.B1(_01705_),
    .VDD(VPWR),
    .Y(_01706_),
    .VSS(VGND),
    .A1(_01495_),
    .A2(_01701_));
 sg13g2_o21ai_1 _07346_ (.B1(_01706_),
    .VDD(VPWR),
    .Y(_01477_),
    .VSS(VGND),
    .A1(\acc_sub.reg2en.q[0] ),
    .A2(_01700_));
 sg13g2_inv_1 _07347_ (.VDD(VPWR),
    .Y(_01707_),
    .A(\acc_sub.add_renorm0.mantisa[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07348_ (.Y(_01708_),
    .A(_01587_),
    .B(\acc_sub.reg2en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07349_ (.B1(_01708_),
    .VDD(VPWR),
    .Y(_01476_),
    .VSS(VGND),
    .A1(\acc_sub.reg2en.q[0] ),
    .A2(_01707_));
 sg13g2_inv_1 _07350_ (.VDD(VPWR),
    .Y(_01709_),
    .A(\acc_sub.add_renorm0.exp[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07351_ (.Y(_01710_),
    .A(net1799),
    .B(\acc_sub.seg_reg0.q[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07352_ (.B1(_01710_),
    .VDD(VPWR),
    .Y(_01475_),
    .VSS(VGND),
    .A1(net1797),
    .A2(_01709_));
 sg13g2_inv_1 _07353_ (.VDD(VPWR),
    .Y(_01711_),
    .A(\acc_sub.add_renorm0.exp[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07354_ (.Y(_01712_),
    .A(net1797),
    .B(\acc_sub.seg_reg0.q[28] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07355_ (.B1(_01712_),
    .VDD(VPWR),
    .Y(_01474_),
    .VSS(VGND),
    .A1(net1797),
    .A2(_01711_));
 sg13g2_inv_2 _07356_ (.Y(_01713_),
    .A(\acc_sub.add_renorm0.exp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07357_ (.Y(_01714_),
    .A(net1799),
    .B(\acc_sub.seg_reg0.q[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07358_ (.B1(_01714_),
    .VDD(VPWR),
    .Y(_01473_),
    .VSS(VGND),
    .A1(net1799),
    .A2(_01713_));
 sg13g2_inv_2 _07359_ (.Y(_01715_),
    .A(\acc_sub.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07360_ (.Y(_01716_),
    .A(net1799),
    .B(\acc_sub.seg_reg0.q[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07361_ (.B1(_01716_),
    .VDD(VPWR),
    .Y(_01472_),
    .VSS(VGND),
    .A1(net1798),
    .A2(_01715_));
 sg13g2_inv_1 _07362_ (.VDD(VPWR),
    .Y(_01717_),
    .A(\acc_sub.add_renorm0.exp[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07363_ (.Y(_01718_),
    .A(net1799),
    .B(\acc_sub.seg_reg0.q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07364_ (.B1(_01718_),
    .VDD(VPWR),
    .Y(_01471_),
    .VSS(VGND),
    .A1(net1798),
    .A2(_01717_));
 sg13g2_inv_1 _07365_ (.VDD(VPWR),
    .Y(_01719_),
    .A(\acc_sub.add_renorm0.exp[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07366_ (.Y(_01720_),
    .A(net1799),
    .B(\acc_sub.seg_reg0.q[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07367_ (.B1(_01720_),
    .VDD(VPWR),
    .Y(_01470_),
    .VSS(VGND),
    .A1(net1798),
    .A2(_01719_));
 sg13g2_inv_2 _07368_ (.Y(_01721_),
    .A(\acc_sub.add_renorm0.exp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07369_ (.Y(_01722_),
    .A(net1799),
    .B(\acc_sub.seg_reg0.q[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07370_ (.B1(_01722_),
    .VDD(VPWR),
    .Y(_01469_),
    .VSS(VGND),
    .A1(net1798),
    .A2(_01721_));
 sg13g2_mux2_1 _07371_ (.A0(\acc_sub.add_renorm0.exp[0] ),
    .A1(\acc_sub.seg_reg0.q[22] ),
    .S(net1797),
    .X(_01468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07372_ (.Y(_01723_),
    .A(\acc[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07373_ (.A(\acc_sub.exp_mant_logic0.a[15] ),
    .B(net1893),
    .Y(_01724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07374_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01723_),
    .A2(net1893),
    .Y(_01467_),
    .B1(_01724_));
 sg13g2_inv_1 _07375_ (.VDD(VPWR),
    .Y(_01725_),
    .A(\acc_sub.exp_mant_logic0.a[14] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07376_ (.Y(_01726_),
    .A(net1886),
    .B(\acc[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07377_ (.B1(_01726_),
    .VDD(VPWR),
    .Y(_01466_),
    .VSS(VGND),
    .A1(net1886),
    .A2(_01725_));
 sg13g2_inv_2 _07378_ (.Y(_01727_),
    .A(\acc_sub.exp_mant_logic0.a[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07379_ (.Y(_01728_),
    .A(net1888),
    .B(\acc[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07380_ (.B1(_01728_),
    .VDD(VPWR),
    .Y(_01465_),
    .VSS(VGND),
    .A1(net1887),
    .A2(_01727_));
 sg13g2_inv_1 _07381_ (.VDD(VPWR),
    .Y(_01729_),
    .A(\acc_sub.exp_mant_logic0.a[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07382_ (.Y(_01730_),
    .A(net1886),
    .B(\acc[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07383_ (.B1(_01730_),
    .VDD(VPWR),
    .Y(_01464_),
    .VSS(VGND),
    .A1(net1886),
    .A2(_01729_));
 sg13g2_inv_2 _07384_ (.Y(_01731_),
    .A(\acc_sub.exp_mant_logic0.a[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07385_ (.Y(_01732_),
    .A(\acc_sub.reg1en.d[0] ),
    .B(\acc[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07386_ (.B1(_01732_),
    .VDD(VPWR),
    .Y(_01463_),
    .VSS(VGND),
    .A1(\acc_sub.reg1en.d[0] ),
    .A2(_01731_));
 sg13g2_inv_1 _07387_ (.VDD(VPWR),
    .Y(_01733_),
    .A(\acc_sub.exp_mant_logic0.a[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07388_ (.Y(_01734_),
    .A(net1893),
    .B(\acc[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07389_ (.B1(_01734_),
    .VDD(VPWR),
    .Y(_01462_),
    .VSS(VGND),
    .A1(net1893),
    .A2(_01733_));
 sg13g2_inv_1 _07390_ (.VDD(VPWR),
    .Y(_01735_),
    .A(\acc_sub.exp_mant_logic0.a[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07391_ (.Y(_01736_),
    .A(net1894),
    .B(\acc[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07392_ (.B1(_01736_),
    .VDD(VPWR),
    .Y(_01461_),
    .VSS(VGND),
    .A1(net1895),
    .A2(_01735_));
 sg13g2_inv_1 _07393_ (.VDD(VPWR),
    .Y(_01737_),
    .A(\acc_sub.exp_mant_logic0.a[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07394_ (.Y(_01738_),
    .A(net1893),
    .B(\acc[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07395_ (.B1(_01738_),
    .VDD(VPWR),
    .Y(_01460_),
    .VSS(VGND),
    .A1(net1895),
    .A2(_01737_));
 sg13g2_inv_2 _07396_ (.Y(_01739_),
    .A(\acc_sub.exp_mant_logic0.a[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07397_ (.Y(_01740_),
    .A(net1893),
    .B(\acc[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07398_ (.B1(_01740_),
    .VDD(VPWR),
    .Y(_01459_),
    .VSS(VGND),
    .A1(net1895),
    .A2(_01739_));
 sg13g2_inv_1 _07399_ (.VDD(VPWR),
    .Y(_01741_),
    .A(\acc_sub.exp_mant_logic0.a[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07400_ (.Y(_01742_),
    .A(net1890),
    .B(\acc[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07401_ (.B1(_01742_),
    .VDD(VPWR),
    .Y(_01458_),
    .VSS(VGND),
    .A1(net1890),
    .A2(_01741_));
 sg13g2_inv_2 _07402_ (.Y(_01743_),
    .A(\acc_sub.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07403_ (.Y(_01744_),
    .A(net1887),
    .B(\acc[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07404_ (.B1(_01744_),
    .VDD(VPWR),
    .Y(_01457_),
    .VSS(VGND),
    .A1(net1890),
    .A2(_01743_));
 sg13g2_inv_2 _07405_ (.Y(_01745_),
    .A(\acc_sub.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07406_ (.Y(_01746_),
    .A(net1894),
    .B(\acc[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07407_ (.B1(_01746_),
    .VDD(VPWR),
    .Y(_01456_),
    .VSS(VGND),
    .A1(net1889),
    .A2(_01745_));
 sg13g2_inv_2 _07408_ (.Y(_01747_),
    .A(\acc_sub.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07409_ (.Y(_01748_),
    .A(net1889),
    .B(\acc[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07410_ (.B1(_01748_),
    .VDD(VPWR),
    .Y(_01455_),
    .VSS(VGND),
    .A1(net1891),
    .A2(_01747_));
 sg13g2_inv_1 _07411_ (.VDD(VPWR),
    .Y(_01749_),
    .A(\acc_sub.exp_mant_logic0.a[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07412_ (.Y(_01750_),
    .A(net1894),
    .B(\acc[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07413_ (.B1(_01750_),
    .VDD(VPWR),
    .Y(_01454_),
    .VSS(VGND),
    .A1(net1889),
    .A2(_01749_));
 sg13g2_inv_2 _07414_ (.Y(_01751_),
    .A(\acc_sub.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07415_ (.Y(_01752_),
    .A(net1894),
    .B(\acc[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07416_ (.B1(_01752_),
    .VDD(VPWR),
    .Y(_01453_),
    .VSS(VGND),
    .A1(net1894),
    .A2(_01751_));
 sg13g2_inv_2 _07417_ (.Y(_01753_),
    .A(\acc_sub.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07418_ (.Y(_01754_),
    .A(net1890),
    .B(\acc[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07419_ (.B1(_01754_),
    .VDD(VPWR),
    .Y(_01452_),
    .VSS(VGND),
    .A1(net1890),
    .A2(_01753_));
 sg13g2_inv_1 _07420_ (.VDD(VPWR),
    .Y(_01755_),
    .A(\fpdiv.reg1en.q[0] ),
    .VSS(VGND));
 sg13g2_nor2_2 _07421_ (.A(\fpdiv.divider0.state ),
    .B(_01755_),
    .Y(_01756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout64 (.A(net67),
    .X(net64),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07423_ (.VDD(VPWR),
    .Y(_01758_),
    .A(_01756_),
    .VSS(VGND));
 sg13g2_inv_1 _07424_ (.VDD(VPWR),
    .Y(_01759_),
    .A(\fpdiv.divider0.divisor_reg[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07425_ (.Y(_01451_),
    .A(_01758_),
    .B(_01759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07426_ (.VDD(VPWR),
    .Y(_01760_),
    .A(\fpdiv.divider0.divisor_reg[10] ),
    .VSS(VGND));
 sg13g2_buf_2 place1775 (.A(net1774),
    .X(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07428_ (.Y(_01762_),
    .A(net1749),
    .B(\fpdiv.divider0.divisor[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07429_ (.B1(_01762_),
    .VDD(VPWR),
    .Y(_01450_),
    .VSS(VGND),
    .A1(_01760_),
    .A2(_01756_));
 sg13g2_inv_1 _07430_ (.VDD(VPWR),
    .Y(_01763_),
    .A(\fpdiv.divider0.divisor[9] ),
    .VSS(VGND));
 sg13g2_buf_2 place1760 (.A(net1759),
    .X(net1760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07432_ (.A(\fpdiv.divider0.divisor_reg[9] ),
    .B(net1749),
    .Y(_01765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07433_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01763_),
    .A2(net1749),
    .Y(_01449_),
    .B1(_01765_));
 sg13g2_inv_1 _07434_ (.VDD(VPWR),
    .Y(_01766_),
    .A(\fpdiv.divider0.divisor[8] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07435_ (.A(\fpdiv.divider0.divisor_reg[8] ),
    .B(net1750),
    .Y(_01767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01766_),
    .A2(net1750),
    .Y(_01448_),
    .B1(_01767_));
 sg13g2_inv_1 _07437_ (.VDD(VPWR),
    .Y(_01768_),
    .A(\fpdiv.divider0.divisor[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07438_ (.A(\fpdiv.divider0.divisor_reg[7] ),
    .B(net1749),
    .Y(_01769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07439_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01768_),
    .A2(net1749),
    .Y(_01447_),
    .B1(_01769_));
 sg13g2_inv_1 _07440_ (.VDD(VPWR),
    .Y(_01770_),
    .A(\fpdiv.divider0.divisor_reg[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07441_ (.Y(_01771_),
    .A(net1749),
    .B(\fpdiv.divider0.divisor[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07442_ (.B1(_01771_),
    .VDD(VPWR),
    .Y(_01446_),
    .VSS(VGND),
    .A1(_01770_),
    .A2(net1750));
 sg13g2_inv_1 _07443_ (.VDD(VPWR),
    .Y(_01772_),
    .A(\fpdiv.divider0.divisor_reg[5] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07444_ (.Y(_01773_),
    .A(net1750),
    .B(\fpdiv.divider0.divisor[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07445_ (.B1(_01773_),
    .VDD(VPWR),
    .Y(_01445_),
    .VSS(VGND),
    .A1(_01772_),
    .A2(net1750));
 sg13g2_inv_1 _07446_ (.VDD(VPWR),
    .Y(_01774_),
    .A(\fpdiv.divider0.divisor_reg[4] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07447_ (.Y(_01775_),
    .A(net1750),
    .B(\fpdiv.divider0.divisor[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07448_ (.B1(_01775_),
    .VDD(VPWR),
    .Y(_01444_),
    .VSS(VGND),
    .A1(_01774_),
    .A2(net1748));
 sg13g2_or2_1 _07449_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_01443_),
    .B(\acc_sub.reg_add_sub.q[0] ),
    .A(net1895));
 sg13g2_mux2_1 _07450_ (.A0(\acc_sub.op_sign_logic0.s_a ),
    .A1(\acc_sub.exp_mant_logic0.a[15] ),
    .S(net1796),
    .X(_01442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07451_ (.Y(_01776_),
    .A(\acc_sub.exp_mant_logic0.b[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07452_ (.A(net1796),
    .B(\acc_sub.op_sign_logic0.s_b ),
    .Y(_01777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07453_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1796),
    .A2(_01776_),
    .Y(_01441_),
    .B1(_01777_));
 sg13g2_mux2_1 _07454_ (.A0(\acc_sub.op_sign_logic0.add_sub ),
    .A1(\acc_sub.reg_add_sub.q[0] ),
    .S(\acc_sub.reg1en.q[0] ),
    .X(_01440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07455_ (.VDD(VPWR),
    .Y(_01778_),
    .A(\acc_sub.seg_reg0.q[29] ),
    .VSS(VGND));
 sg13g2_inv_4 _07456_ (.A(\acc_sub.reg1en.q[0] ),
    .Y(_01779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout48 (.A(net49),
    .X(net48),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout46 (.A(net47),
    .X(net46),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07459_ (.A(\acc_sub.exp_mant_logic0.b[14] ),
    .B(net1782),
    .Y(_01782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07460_ (.A(\acc_sub.exp_mant_logic0.b[13] ),
    .B(_01727_),
    .Y(_01783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07461_ (.VDD(VPWR),
    .Y(_01784_),
    .A(\acc_sub.exp_mant_logic0.b[13] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07462_ (.A(\acc_sub.exp_mant_logic0.a[13] ),
    .B(_01784_),
    .Y(_01785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07463_ (.A(_01783_),
    .B(_01785_),
    .Y(_01786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07464_ (.VDD(VPWR),
    .Y(_01787_),
    .A(_01786_),
    .VSS(VGND));
 sg13g2_nor2_1 _07465_ (.A(\acc_sub.exp_mant_logic0.b[14] ),
    .B(_01725_),
    .Y(_01788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07466_ (.VDD(VPWR),
    .Y(_01789_),
    .A(\acc_sub.exp_mant_logic0.b[14] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07467_ (.A(\acc_sub.exp_mant_logic0.a[14] ),
    .B(_01789_),
    .Y(_01790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07468_ (.A(_01788_),
    .B(_01790_),
    .Y(_01791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07469_ (.VDD(VPWR),
    .Y(_01792_),
    .A(_01791_),
    .VSS(VGND));
 sg13g2_nor2_1 _07470_ (.A(_01787_),
    .B(_01792_),
    .Y(_01793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07471_ (.A(\acc_sub.exp_mant_logic0.b[12] ),
    .B(_01729_),
    .Y(_01794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07472_ (.VDD(VPWR),
    .Y(_01795_),
    .A(\acc_sub.exp_mant_logic0.b[12] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07473_ (.A(\acc_sub.exp_mant_logic0.a[12] ),
    .B(_01795_),
    .Y(_01796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07474_ (.A(_01794_),
    .B(_01796_),
    .Y(_01797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07475_ (.A(\acc_sub.exp_mant_logic0.b[11] ),
    .B(_01731_),
    .Y(_01798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07476_ (.VDD(VPWR),
    .Y(_01799_),
    .A(\acc_sub.exp_mant_logic0.b[11] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07477_ (.A(\acc_sub.exp_mant_logic0.a[11] ),
    .B(_01799_),
    .Y(_01800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07478_ (.A(_01798_),
    .B(_01800_),
    .Y(_01801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _07479_ (.X(_01802_),
    .A(_01793_),
    .B(_01797_),
    .C(_01801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07480_ (.A(\acc_sub.exp_mant_logic0.b[10] ),
    .B(_01733_),
    .Y(_01803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07481_ (.Y(_01804_),
    .A(\acc_sub.exp_mant_logic0.b[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07482_ (.A(\acc_sub.exp_mant_logic0.a[10] ),
    .B(_01804_),
    .Y(_01805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07483_ (.A(_01803_),
    .B(_01805_),
    .Y(_01806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07484_ (.A(\acc_sub.exp_mant_logic0.b[9] ),
    .B(_01735_),
    .Y(_01807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07485_ (.VDD(VPWR),
    .Y(_01808_),
    .A(\acc_sub.exp_mant_logic0.b[9] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07486_ (.A(\acc_sub.exp_mant_logic0.a[9] ),
    .B(_01808_),
    .Y(_01809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07487_ (.A(_01807_),
    .B(_01809_),
    .Y(_01810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07488_ (.Y(_01811_),
    .A(_01806_),
    .B(_01810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _07489_ (.B(\acc_sub.exp_mant_logic0.b[8] ),
    .A(\acc_sub.exp_mant_logic0.a[8] ),
    .X(_01812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07490_ (.VDD(VPWR),
    .Y(_01813_),
    .A(\acc_sub.exp_mant_logic0.b[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07491_ (.A(\acc_sub.exp_mant_logic0.a[7] ),
    .B(_01813_),
    .Y(_01814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07492_ (.A(\acc_sub.exp_mant_logic0.b[7] ),
    .B(_01739_),
    .Y(_01815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07493_ (.A(_01814_),
    .B(_01815_),
    .Y(_01816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07494_ (.VDD(VPWR),
    .Y(_01817_),
    .A(_01816_),
    .VSS(VGND));
 sg13g2_nor2_1 _07495_ (.A(_01812_),
    .B(_01817_),
    .Y(_01818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07496_ (.VDD(VPWR),
    .Y(_01819_),
    .A(_01818_),
    .VSS(VGND));
 sg13g2_nor2_1 _07497_ (.A(_01811_),
    .B(_01819_),
    .Y(_01820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07498_ (.Y(_01821_),
    .A(_01802_),
    .B(_01820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1709 (.A(_04775_),
    .X(net1709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07500_ (.Y(_01823_),
    .A(_01821_),
    .B(\acc_sub.exp_mant_logic0.a[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07501_ (.Y(_01439_),
    .B1(_01782_),
    .B2(_01823_),
    .A2(net1782),
    .A1(_01778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07502_ (.VDD(VPWR),
    .Y(_01824_),
    .A(\acc_sub.seg_reg0.q[28] ),
    .VSS(VGND));
 sg13g2_inv_1 _07503_ (.VDD(VPWR),
    .Y(_01825_),
    .A(\acc_sub.exp_mant_logic0.b[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07504_ (.Y(_01826_),
    .A(_01825_),
    .B(\acc_sub.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07505_ (.B1(_01826_),
    .VDD(VPWR),
    .Y(_01827_),
    .VSS(VGND),
    .A1(_01814_),
    .A2(_01812_));
 sg13g2_nand2_1 _07506_ (.Y(_01828_),
    .A(_01827_),
    .B(_01810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07507_ (.Y(_01829_),
    .B(_01828_),
    .A_N(_01807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07508_ (.VDD(VPWR),
    .Y(_01830_),
    .A(_01805_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07509_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01829_),
    .A2(_01830_),
    .Y(_01831_),
    .B1(_01803_));
 sg13g2_inv_1 _07510_ (.VDD(VPWR),
    .Y(_01832_),
    .A(_01831_),
    .VSS(VGND));
 sg13g2_nand2_1 _07511_ (.Y(_01833_),
    .A(_01832_),
    .B(_01802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07512_ (.VDD(VPWR),
    .Y(_01834_),
    .A(_01796_),
    .VSS(VGND));
 sg13g2_a21o_1 _07513_ (.A2(_01798_),
    .A1(_01834_),
    .B1(_01794_),
    .X(_01835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _07514_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_01793_),
    .C1(_01788_),
    .B1(_01835_),
    .A1(_01783_),
    .Y(_01836_),
    .A2(_01791_));
 sg13g2_nand2_2 _07515_ (.Y(_01837_),
    .A(_01833_),
    .B(_01836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07516_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01837_),
    .A2(_01727_),
    .Y(_01838_),
    .B1(net1782));
 sg13g2_o21ai_1 _07517_ (.B1(_01838_),
    .VDD(VPWR),
    .Y(_01839_),
    .VSS(VGND),
    .A1(\acc_sub.exp_mant_logic0.b[13] ),
    .A2(_01837_));
 sg13g2_o21ai_1 _07518_ (.B1(_01839_),
    .VDD(VPWR),
    .Y(_01438_),
    .VSS(VGND),
    .A1(_01824_),
    .A2(net1796));
 sg13g2_nand2_1 _07519_ (.Y(_01840_),
    .A(_01837_),
    .B(_01821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07522_ (.VDD(VPWR),
    .Y(_01843_),
    .A(net1686),
    .VSS(VGND));
 sg13g2_nor2_2 _07523_ (.A(_01779_),
    .B(_01843_),
    .Y(_01844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07525_ (.Y(_01846_),
    .A(_01844_),
    .B(\acc_sub.exp_mant_logic0.b[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07526_ (.A(net1782),
    .B(_01840_),
    .Y(_01847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07529_ (.Y(_01850_),
    .A(_01847_),
    .B(\acc_sub.exp_mant_logic0.a[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07530_ (.Y(_01851_),
    .A(net1782),
    .B(\acc_sub.seg_reg0.q[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07531_ (.B(_01850_),
    .C(_01851_),
    .A(_01846_),
    .Y(_01437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07532_ (.Y(_01852_),
    .A(_01844_),
    .B(\acc_sub.exp_mant_logic0.b[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07533_ (.Y(_01853_),
    .A(_01847_),
    .B(\acc_sub.exp_mant_logic0.a[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07534_ (.Y(_01854_),
    .A(net1782),
    .B(\acc_sub.seg_reg0.q[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07535_ (.B(_01853_),
    .C(_01854_),
    .A(_01852_),
    .Y(_01436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07536_ (.Y(_01855_),
    .A(_01844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07537_ (.Y(_01856_),
    .B1(\acc_sub.exp_mant_logic0.a[10] ),
    .B2(_01847_),
    .A2(_01779_),
    .A1(\acc_sub.seg_reg0.q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07538_ (.B1(_01856_),
    .VDD(VPWR),
    .Y(_01435_),
    .VSS(VGND),
    .A1(_01804_),
    .A2(_01855_));
 sg13g2_nand2_1 _07539_ (.Y(_01857_),
    .A(_01844_),
    .B(\acc_sub.exp_mant_logic0.b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07540_ (.Y(_01858_),
    .A(_01847_),
    .B(\acc_sub.exp_mant_logic0.a[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07541_ (.Y(_01859_),
    .A(_01779_),
    .B(\acc_sub.seg_reg0.q[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07542_ (.B(_01858_),
    .C(_01859_),
    .A(_01857_),
    .Y(_01434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07543_ (.Y(_01860_),
    .A(_01844_),
    .B(\acc_sub.exp_mant_logic0.b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07544_ (.Y(_01861_),
    .A(_01847_),
    .B(\acc_sub.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07545_ (.Y(_01862_),
    .A(_01779_),
    .B(\acc_sub.seg_reg0.q[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07546_ (.B(_01861_),
    .C(_01862_),
    .A(_01860_),
    .Y(_01433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07547_ (.Y(_01863_),
    .B1(\acc_sub.exp_mant_logic0.a[7] ),
    .B2(_01847_),
    .A2(_01779_),
    .A1(\acc_sub.seg_reg0.q[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07548_ (.B1(_01863_),
    .VDD(VPWR),
    .Y(_01432_),
    .VSS(VGND),
    .A1(_01813_),
    .A2(_01855_));
 sg13g2_nand3_1 _07549_ (.B(_01745_),
    .C(_01751_),
    .A(_01743_),
    .Y(_01864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _07550_ (.B(_01735_),
    .C(_01737_),
    .A(_01733_),
    .Y(_01865_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01739_));
 sg13g2_nand4_1 _07551_ (.B(_01727_),
    .C(_01729_),
    .A(_01725_),
    .Y(_01866_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01731_));
 sg13g2_nand4_1 _07552_ (.B(_01747_),
    .C(_01749_),
    .A(_01741_),
    .Y(_01867_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_01753_));
 sg13g2_nor4_2 _07553_ (.A(_01864_),
    .B(_01865_),
    .C(_01866_),
    .Y(_01868_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01867_));
 sg13g2_inv_4 _07554_ (.A(_01868_),
    .Y(_01869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07555_ (.B(net1796),
    .C(_01869_),
    .A(_01837_),
    .Y(_01870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07556_ (.B1(_01870_),
    .VDD(VPWR),
    .Y(_01431_),
    .VSS(VGND),
    .A1(\acc_sub.reg1en.q[0] ),
    .A2(_01499_));
 sg13g2_inv_4 _07557_ (.A(_01821_),
    .Y(_01871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1691 (.A(_02275_),
    .X(net1691),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07559_ (.VDD(VPWR),
    .Y(_01873_),
    .A(_01801_),
    .VSS(VGND));
 sg13g2_inv_1 _07560_ (.VDD(VPWR),
    .Y(_01874_),
    .A(_01798_),
    .VSS(VGND));
 sg13g2_o21ai_1 _07561_ (.B1(_01874_),
    .VDD(VPWR),
    .Y(_01875_),
    .VSS(VGND),
    .A1(_01873_),
    .A2(_01831_));
 sg13g2_a21oi_1 _07562_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01875_),
    .A2(_01834_),
    .Y(_01876_),
    .B1(_01794_));
 sg13g2_inv_1 _07563_ (.VDD(VPWR),
    .Y(_01877_),
    .A(_01783_),
    .VSS(VGND));
 sg13g2_o21ai_1 _07564_ (.B1(_01877_),
    .VDD(VPWR),
    .Y(_01878_),
    .VSS(VGND),
    .A1(_01787_),
    .A2(_01876_));
 sg13g2_nand2b_1 _07565_ (.Y(_01879_),
    .B(_01878_),
    .A_N(_01790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07566_ (.VDD(VPWR),
    .Y(_01880_),
    .A(_01812_),
    .VSS(VGND));
 sg13g2_inv_1 _07567_ (.VDD(VPWR),
    .Y(_01881_),
    .A(_01815_),
    .VSS(VGND));
 sg13g2_nand2_1 _07568_ (.Y(_01882_),
    .A(_01880_),
    .B(_01881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07569_ (.B1(_01882_),
    .VDD(VPWR),
    .Y(_01883_),
    .VSS(VGND),
    .A1(\acc_sub.exp_mant_logic0.a[8] ),
    .A2(_01825_));
 sg13g2_inv_1 _07570_ (.VDD(VPWR),
    .Y(_01884_),
    .A(_01883_),
    .VSS(VGND));
 sg13g2_nor2_1 _07571_ (.A(_01811_),
    .B(_01884_),
    .Y(_01885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07572_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01806_),
    .A2(_01809_),
    .Y(_01886_),
    .B1(_01805_));
 sg13g2_nor2b_1 _07573_ (.A(_01885_),
    .B_N(_01886_),
    .Y(_01887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07574_ (.VDD(VPWR),
    .Y(_01888_),
    .A(_01887_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07575_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01888_),
    .A2(_01801_),
    .Y(_01889_),
    .B1(_01800_));
 sg13g2_o21ai_1 _07576_ (.B1(_01834_),
    .VDD(VPWR),
    .Y(_01890_),
    .VSS(VGND),
    .A1(_01794_),
    .A2(_01889_));
 sg13g2_a21oi_1 _07577_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01890_),
    .A2(_01786_),
    .Y(_01891_),
    .B1(_01785_));
 sg13g2_nand2b_1 _07578_ (.Y(_01892_),
    .B(net1687),
    .A_N(_01891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07579_ (.B1(_01892_),
    .VDD(VPWR),
    .Y(_01893_),
    .VSS(VGND),
    .A1(_01871_),
    .A2(_01879_));
 sg13g2_nand2_1 _07580_ (.Y(_01894_),
    .A(_01890_),
    .B(net1687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07581_ (.B1(_01894_),
    .VDD(VPWR),
    .Y(_01895_),
    .VSS(VGND),
    .A1(net1687),
    .A2(_01876_));
 sg13g2_xnor2_1 _07582_ (.Y(_01896_),
    .A(_01787_),
    .B(_01895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07583_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01893_),
    .A2(_01792_),
    .Y(_01897_),
    .B1(_01896_));
 sg13g2_nand2_1 _07584_ (.Y(_01898_),
    .A(net1687),
    .B(_01889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07585_ (.B1(_01898_),
    .VDD(VPWR),
    .Y(_01899_),
    .VSS(VGND),
    .A1(_01875_),
    .A2(net1687));
 sg13g2_xnor2_1 _07586_ (.Y(_01900_),
    .A(_01797_),
    .B(_01899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07587_ (.A(_01832_),
    .B(net1687),
    .Y(_01901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07588_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1687),
    .A2(_01887_),
    .Y(_01902_),
    .B1(_01901_));
 sg13g2_xnor2_1 _07589_ (.Y(_01903_),
    .A(_01873_),
    .B(_01902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07590_ (.A(_01900_),
    .B(_01903_),
    .Y(_01904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07591_ (.Y(_01905_),
    .A(_01897_),
    .B(_01904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07592_ (.Y(_01906_),
    .A(net1686),
    .B(_01881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07593_ (.B1(_01906_),
    .VDD(VPWR),
    .Y(_01907_),
    .VSS(VGND),
    .A1(_01814_),
    .A2(net1686));
 sg13g2_xnor2_1 _07594_ (.Y(_01908_),
    .A(_01812_),
    .B(_01907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07595_ (.VDD(VPWR),
    .Y(_01909_),
    .A(_01908_),
    .VSS(VGND));
 sg13g2_nand2_1 _07596_ (.Y(_01910_),
    .A(_01909_),
    .B(_01817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07597_ (.Y(_01911_),
    .A(net1686),
    .B(_01884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07598_ (.B1(_01911_),
    .VDD(VPWR),
    .Y(_01912_),
    .VSS(VGND),
    .A1(_01827_),
    .A2(net1686));
 sg13g2_xor2_1 _07599_ (.B(_01912_),
    .A(_01810_),
    .X(_01913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07600_ (.VDD(VPWR),
    .Y(_01914_),
    .A(_01913_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07601_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01883_),
    .A2(_01810_),
    .Y(_01915_),
    .B1(_01809_));
 sg13g2_nor2_1 _07602_ (.A(_01829_),
    .B(net1686),
    .Y(_01916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1686),
    .A2(_01915_),
    .Y(_01917_),
    .B1(_01916_));
 sg13g2_xnor2_1 _07604_ (.Y(_01918_),
    .A(_01806_),
    .B(_01917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07605_ (.VDD(VPWR),
    .Y(_01919_),
    .A(_01918_),
    .VSS(VGND));
 sg13g2_nor2_1 _07606_ (.A(_01914_),
    .B(_01919_),
    .Y(_01920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07607_ (.VDD(VPWR),
    .Y(_01921_),
    .A(_01920_),
    .VSS(VGND));
 sg13g2_nor2_1 _07608_ (.A(_01910_),
    .B(_01921_),
    .Y(_01922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _07609_ (.A(net1660),
    .B_N(_01922_),
    .Y(_01923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_83_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_83_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_82_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_82_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07612_ (.Y(_01926_),
    .B1(_01869_),
    .B2(_01923_),
    .A2(_01871_),
    .A1(net1792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07613_ (.B(_01818_),
    .C(_01913_),
    .A(_01919_),
    .Y(_01927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07614_ (.A(_01816_),
    .B(_01909_),
    .Y(_01928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07615_ (.Y(_01929_),
    .A(_01920_),
    .B(_01928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_54_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_54_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01927_),
    .A2(_01929_),
    .Y(_01931_),
    .B1(net1660));
 sg13g2_nor3_1 _07618_ (.A(_01871_),
    .B(_01923_),
    .C(_01931_),
    .Y(_01932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07619_ (.Y(_01933_),
    .A(_01914_),
    .B(_01918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07620_ (.A(_01819_),
    .B(_01933_),
    .Y(_01934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _07621_ (.A(_01905_),
    .B_N(_01934_),
    .Y(_01935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07622_ (.A(_01880_),
    .B(_01817_),
    .Y(_01936_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07623_ (.VDD(VPWR),
    .Y(_01937_),
    .A(_01936_),
    .VSS(VGND));
 sg13g2_nor2_1 _07624_ (.A(_01937_),
    .B(_01921_),
    .Y(_01938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07625_ (.VDD(VPWR),
    .Y(_01939_),
    .A(_01938_),
    .VSS(VGND));
 sg13g2_inv_1 _07626_ (.VDD(VPWR),
    .Y(_01940_),
    .A(_01933_),
    .VSS(VGND));
 sg13g2_nand2_1 _07627_ (.Y(_01941_),
    .A(_01940_),
    .B(_01819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01939_),
    .A2(_01941_),
    .Y(_01942_),
    .B1(_01905_));
 sg13g2_nor2_1 _07629_ (.A(_01935_),
    .B(_01942_),
    .Y(_01943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01932_),
    .A2(_01943_),
    .Y(_01944_),
    .B1(_01855_));
 sg13g2_buf_8 clkbuf_leaf_95_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_95_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07632_ (.Y(_01946_),
    .B(net1641),
    .A_N(_01926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout45 (.A(net46),
    .X(net45),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07634_ (.Y(_01948_),
    .B1(net1792),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[9] ),
    .A1(net1779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07635_ (.Y(_01430_),
    .A(_01946_),
    .B(_01948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07636_ (.A(_01939_),
    .B(_01905_),
    .Y(_01949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_94_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_94_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_93_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_93_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07639_ (.Y(_01952_),
    .A(net1646),
    .B(_01869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07640_ (.Y(_01953_),
    .A(_01923_),
    .B(net1792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07641_ (.Y(_01954_),
    .A(net1685),
    .B(net1793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07642_ (.B(_01953_),
    .C(_01954_),
    .A(_01952_),
    .Y(_01955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07643_ (.Y(_01956_),
    .A(net1641),
    .B(_01955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07644_ (.Y(_01957_),
    .B1(net1793),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[8] ),
    .A1(net1780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07645_ (.Y(_01429_),
    .A(_01956_),
    .B(_01957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07646_ (.Y(_01958_),
    .B1(net1792),
    .B2(net1646),
    .A2(net1793),
    .A1(net1651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07647_ (.A(_01929_),
    .B(net1660),
    .Y(_01959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_86_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_86_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_85_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_85_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07650_ (.Y(_01962_),
    .B1(_01869_),
    .B2(net1649),
    .A2(net1685),
    .A1(\acc_sub.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07651_ (.Y(_01963_),
    .A(_01958_),
    .B(_01962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07652_ (.Y(_01964_),
    .A(net1641),
    .B(_01963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07653_ (.Y(_01965_),
    .B1(\acc_sub.exp_mant_logic0.a[4] ),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[7] ),
    .A1(net1780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07654_ (.Y(_01428_),
    .A(_01964_),
    .B(_01965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_84_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_84_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07656_ (.Y(_01967_),
    .B1(net1793),
    .B2(net1646),
    .A2(_01869_),
    .A1(_01935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07657_ (.Y(_01968_),
    .A(net1649),
    .B(net1792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07658_ (.Y(_01969_),
    .B1(\acc_sub.exp_mant_logic0.a[4] ),
    .B2(net1651),
    .A2(net1685),
    .A1(\acc_sub.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07659_ (.B(_01968_),
    .C(_01969_),
    .A(_01967_),
    .Y(_01970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07660_ (.Y(_01971_),
    .A(_01970_),
    .B(net1641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07661_ (.Y(_01972_),
    .B1(\acc_sub.exp_mant_logic0.a[3] ),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[6] ),
    .A1(net1780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07662_ (.Y(_01427_),
    .A(_01971_),
    .B(_01972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07663_ (.A(_01749_),
    .B(_01821_),
    .Y(_01973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07664_ (.A(_01910_),
    .B(_01933_),
    .Y(_01974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _07665_ (.A(net1660),
    .B_N(_01974_),
    .Y(_01975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1653 (.A(_05181_),
    .X(net1653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07667_ (.Y(_01977_),
    .A(_01975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07668_ (.A(_01868_),
    .B(_01977_),
    .Y(_01978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07669_ (.Y(_01979_),
    .A(_01923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07670_ (.A(_01747_),
    .B(_01979_),
    .Y(_01980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07671_ (.A(_01973_),
    .B(_01978_),
    .C(_01980_),
    .Y(_01981_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07672_ (.Y(_01982_),
    .A(_01935_),
    .B(net1792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07673_ (.Y(_01983_),
    .B1(net1793),
    .B2(net1649),
    .A2(\acc_sub.exp_mant_logic0.a[4] ),
    .A1(_01949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07674_ (.B(_01982_),
    .C(_01983_),
    .A(_01981_),
    .Y(_01984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07675_ (.Y(_01985_),
    .A(_01984_),
    .B(net1641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07676_ (.Y(_01986_),
    .B1(\acc_sub.exp_mant_logic0.a[2] ),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[5] ),
    .A1(net1780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07677_ (.Y(_01426_),
    .A(_01985_),
    .B(_01986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07678_ (.Y(_01987_),
    .A(_01949_),
    .B(\acc_sub.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07679_ (.A(_01937_),
    .B(_01933_),
    .Y(_01988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _07680_ (.A(net1660),
    .B_N(_01988_),
    .Y(_01989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_87_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_87_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07682_ (.Y(_01991_),
    .A(_01989_),
    .B(_01869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07683_ (.Y(_01992_),
    .A(_01987_),
    .B(_01991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07684_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1793),
    .A2(_01935_),
    .Y(_01993_),
    .B1(_01992_));
 sg13g2_a22oi_1 _07685_ (.Y(_01994_),
    .B1(\acc_sub.exp_mant_logic0.a[2] ),
    .B2(_01923_),
    .A2(_01871_),
    .A1(\acc_sub.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07686_ (.Y(_01995_),
    .B1(\acc_sub.exp_mant_logic0.a[4] ),
    .B2(net1649),
    .A2(net1792),
    .A1(_01975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07687_ (.B(_01994_),
    .C(_01995_),
    .A(_01993_),
    .Y(_01996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07688_ (.Y(_01997_),
    .A(_01996_),
    .B(net1641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07689_ (.Y(_01998_),
    .B1(\acc_sub.exp_mant_logic0.a[1] ),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[4] ),
    .A1(net1780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07690_ (.Y(_01425_),
    .A(_01997_),
    .B(_01998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07691_ (.Y(_01999_),
    .A(_01949_),
    .B(\acc_sub.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07692_ (.Y(_02000_),
    .A(_01989_),
    .B(net1792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07693_ (.Y(_02001_),
    .A(_01935_),
    .B(\acc_sub.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07694_ (.B(_02000_),
    .C(_02001_),
    .A(_01999_),
    .Y(_02002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07695_ (.Y(_02003_),
    .B1(net1793),
    .B2(_01975_),
    .A2(_01871_),
    .A1(\acc_sub.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _07696_ (.A(_02002_),
    .B_N(_02003_),
    .Y(_02004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07697_ (.Y(_02005_),
    .A(_01940_),
    .B(_01928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07698_ (.A(_02005_),
    .B(net1660),
    .Y(_02006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_88_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_88_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07700_ (.Y(_02008_),
    .A(_01959_),
    .B(\acc_sub.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07701_ (.B1(_02008_),
    .VDD(VPWR),
    .Y(_02009_),
    .VSS(VGND),
    .A1(_01751_),
    .A2(_01979_));
 sg13g2_a21oi_1 _07702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01869_),
    .A2(_02006_),
    .Y(_02010_),
    .B1(_02009_));
 sg13g2_nand2_1 _07703_ (.Y(_02011_),
    .A(_02004_),
    .B(_02010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07704_ (.Y(_02012_),
    .A(_02011_),
    .B(_01944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07705_ (.Y(_02013_),
    .B1(\acc_sub.exp_mant_logic0.a[0] ),
    .B2(net1672),
    .A2(\acc_sub.op_sign_logic0.mantisa_a[3] ),
    .A1(net1779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07706_ (.Y(_01424_),
    .A(_02012_),
    .B(_02013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07707_ (.A(_01745_),
    .B(_01977_),
    .Y(_02014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07708_ (.Y(_02015_),
    .A(_01989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07709_ (.A(_01743_),
    .B(_02015_),
    .Y(_02016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07710_ (.Y(_02017_),
    .A(_02006_),
    .B(\acc_sub.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07711_ (.A(_01927_),
    .B(net1660),
    .Y(_02018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07712_ (.Y(_02019_),
    .A(_02018_),
    .B(_01869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07713_ (.Y(_02020_),
    .A(_02017_),
    .B(_02019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07714_ (.A(_02014_),
    .B(_02016_),
    .C(_02020_),
    .Y(_02021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07715_ (.Y(_02022_),
    .A(_01949_),
    .B(\acc_sub.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07716_ (.B1(_02022_),
    .VDD(VPWR),
    .Y(_02023_),
    .VSS(VGND),
    .A1(_01753_),
    .A2(_01979_));
 sg13g2_inv_2 _07717_ (.Y(_02024_),
    .A(net1650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07718_ (.Y(_02025_),
    .A(_01959_),
    .B(\acc_sub.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07719_ (.B1(_02025_),
    .VDD(VPWR),
    .Y(_02026_),
    .VSS(VGND),
    .A1(_01747_),
    .A2(_02024_));
 sg13g2_nor2_1 _07720_ (.A(_02023_),
    .B(_02026_),
    .Y(_02027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07721_ (.Y(_02028_),
    .A(_02021_),
    .B(_02027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07722_ (.Y(_02029_),
    .A(_02028_),
    .B(_01944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07723_ (.Y(_02030_),
    .A(net1780),
    .B(\acc_sub.op_sign_logic0.mantisa_a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07724_ (.Y(_01423_),
    .A(_02029_),
    .B(_02030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07725_ (.Y(_02031_),
    .A(_01959_),
    .B(\acc_sub.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07726_ (.B1(_02031_),
    .VDD(VPWR),
    .Y(_02032_),
    .VSS(VGND),
    .A1(_01745_),
    .A2(_02015_));
 sg13g2_nor2_1 _07727_ (.A(_01747_),
    .B(_01977_),
    .Y(_02033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07728_ (.Y(_02034_),
    .A(_02018_),
    .B(\acc_sub.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07729_ (.Y(_02035_),
    .A(_02006_),
    .B(\acc_sub.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07730_ (.Y(_02036_),
    .A(_02034_),
    .B(_02035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07731_ (.A(_02033_),
    .B(_02036_),
    .Y(_02037_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07732_ (.Y(_02038_),
    .B1(\acc_sub.exp_mant_logic0.a[0] ),
    .B2(_01949_),
    .A2(\acc_sub.exp_mant_logic0.a[2] ),
    .A1(_01935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _07733_ (.B(_02037_),
    .C(_02038_),
    .Y(_02039_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_02032_));
 sg13g2_nand2_1 _07734_ (.Y(_02040_),
    .A(_02039_),
    .B(net1641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07735_ (.Y(_02041_),
    .A(net1779),
    .B(\acc_sub.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07736_ (.Y(_01422_),
    .A(_02040_),
    .B(_02041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07737_ (.VDD(VPWR),
    .Y(_02042_),
    .A(\acc_sub.op_sign_logic0.mantisa_a[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07738_ (.Y(_02043_),
    .A(_02006_),
    .B(\acc_sub.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07739_ (.Y(_02044_),
    .A(_02018_),
    .B(net1793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07740_ (.Y(_02045_),
    .A(_02043_),
    .B(_02044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07741_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc_sub.exp_mant_logic0.a[2] ),
    .A2(_01975_),
    .Y(_02046_),
    .B1(_02045_));
 sg13g2_nor2_1 _07742_ (.A(_01747_),
    .B(_02015_),
    .Y(_02047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07743_ (.VDD(VPWR),
    .Y(_02048_),
    .A(_01959_),
    .VSS(VGND));
 sg13g2_nor2_1 _07744_ (.A(_01753_),
    .B(_02048_),
    .Y(_02049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07745_ (.A(_01751_),
    .B(_02024_),
    .Y(_02050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07746_ (.A(_02047_),
    .B(_02049_),
    .C(_02050_),
    .Y(_02051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07747_ (.Y(_02052_),
    .A(_02046_),
    .B(_02051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07748_ (.Y(_02053_),
    .A(_02052_),
    .B(_01944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07749_ (.B1(_02053_),
    .VDD(VPWR),
    .Y(_01421_),
    .VSS(VGND),
    .A1(net1796),
    .A2(_02042_));
 sg13g2_nor4_1 _07750_ (.A(\acc_sub.exp_mant_logic0.b[10] ),
    .B(\acc_sub.exp_mant_logic0.b[9] ),
    .C(\acc_sub.exp_mant_logic0.b[8] ),
    .D(\acc_sub.exp_mant_logic0.b[7] ),
    .Y(_02054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _07751_ (.A(\acc_sub.exp_mant_logic0.b[14] ),
    .B(\acc_sub.exp_mant_logic0.b[13] ),
    .C(\acc_sub.exp_mant_logic0.b[12] ),
    .D(\acc_sub.exp_mant_logic0.b[11] ),
    .Y(_02055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _07752_ (.A(\acc_sub.exp_mant_logic0.b[6] ),
    .B(\acc_sub.exp_mant_logic0.b[5] ),
    .C(\acc_sub.exp_mant_logic0.b[4] ),
    .D(\acc_sub.exp_mant_logic0.b[3] ),
    .Y(_02056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07753_ (.A(\acc_sub.exp_mant_logic0.b[2] ),
    .B(\acc_sub.exp_mant_logic0.b[1] ),
    .C(\acc_sub.exp_mant_logic0.b[0] ),
    .Y(_02057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _07754_ (.B(_02055_),
    .C(_02056_),
    .A(_02054_),
    .Y(_02058_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02057_));
 sg13g2_buf_2 place1776 (.A(net1775),
    .X(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07756_ (.B(net1796),
    .C(_02058_),
    .A(net1686),
    .Y(_02060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07757_ (.B1(_02060_),
    .VDD(VPWR),
    .Y(_01420_),
    .VSS(VGND),
    .A1(\acc_sub.reg1en.q[0] ),
    .A2(_01501_));
 sg13g2_a22oi_1 _07758_ (.Y(_02061_),
    .B1(net1747),
    .B2(net1651),
    .A2(net1685),
    .A1(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07759_ (.VDD(VPWR),
    .Y(_02062_),
    .A(_01847_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07760_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01932_),
    .A2(_01943_),
    .Y(_02063_),
    .B1(_02062_));
 sg13g2_buf_8 clkbuf_leaf_96_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_96_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _07762_ (.Y(_02065_),
    .B(net1640),
    .A_N(_02061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07763_ (.Y(_02066_),
    .B1(net1794),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[9] ),
    .A1(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07764_ (.Y(_01419_),
    .A(_02065_),
    .B(_02066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07765_ (.Y(_02067_),
    .A(net1646),
    .B(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07766_ (.Y(_02068_),
    .A(net1651),
    .B(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07767_ (.Y(_02069_),
    .A(net1685),
    .B(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07768_ (.B(_02068_),
    .C(_02069_),
    .A(_02067_),
    .Y(_02070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07769_ (.Y(_02071_),
    .A(net1640),
    .B(_02070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07770_ (.Y(_02072_),
    .B1(net1795),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[8] ),
    .A1(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07771_ (.Y(_01418_),
    .A(_02071_),
    .B(_02072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07772_ (.Y(_02073_),
    .A(\acc_sub.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07773_ (.A(_02073_),
    .B(_01821_),
    .Y(_02074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07774_ (.Y(_02075_),
    .A(net1646),
    .B(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07775_ (.Y(_02076_),
    .A(net1649),
    .B(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07776_ (.Y(_02077_),
    .A(net1651),
    .B(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07777_ (.B(_02076_),
    .C(_02077_),
    .A(_02075_),
    .Y(_02078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07778_ (.B1(net1640),
    .VDD(VPWR),
    .Y(_02079_),
    .VSS(VGND),
    .A1(_02074_),
    .A2(_02078_));
 sg13g2_a22oi_1 _07779_ (.Y(_02080_),
    .B1(\acc_sub.exp_mant_logic0.b[4] ),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[7] ),
    .A1(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07780_ (.Y(_01417_),
    .A(_02079_),
    .B(_02080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07781_ (.Y(_02081_),
    .B1(net1795),
    .B2(net1646),
    .A2(net1747),
    .A1(net1650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07782_ (.Y(_02082_),
    .A(net1649),
    .B(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07783_ (.Y(_02083_),
    .B1(\acc_sub.exp_mant_logic0.b[4] ),
    .B2(net1651),
    .A2(net1685),
    .A1(\acc_sub.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07784_ (.B(_02082_),
    .C(_02083_),
    .A(_02081_),
    .Y(_02084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07785_ (.Y(_02085_),
    .A(_02084_),
    .B(net1640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07786_ (.Y(_02086_),
    .B1(\acc_sub.exp_mant_logic0.b[3] ),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[6] ),
    .A1(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07787_ (.Y(_01416_),
    .A(_02085_),
    .B(_02086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07788_ (.VDD(VPWR),
    .Y(_02087_),
    .A(\acc_sub.exp_mant_logic0.b[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07789_ (.A(_02087_),
    .B(_01821_),
    .Y(_02088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07790_ (.Y(_02089_),
    .A(\acc_sub.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07791_ (.A(_02089_),
    .B(_01979_),
    .Y(_02090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07792_ (.VDD(VPWR),
    .Y(_02091_),
    .A(\acc_sub.exp_mant_logic0.b[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07793_ (.A(_02091_),
    .B(_02048_),
    .Y(_02092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07794_ (.A(_02088_),
    .B(_02090_),
    .C(_02092_),
    .Y(_02093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07795_ (.Y(_02094_),
    .A(_01975_),
    .B(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07796_ (.A(_02073_),
    .B(_01939_),
    .C(_01905_),
    .Y(_02095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07797_ (.VDD(VPWR),
    .Y(_02096_),
    .A(\acc_sub.exp_mant_logic0.b[6] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07798_ (.A(_02096_),
    .B(_02024_),
    .Y(_02097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07799_ (.A(_02095_),
    .B(_02097_),
    .Y(_02098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07800_ (.B(_02094_),
    .C(_02098_),
    .A(_02093_),
    .Y(_02099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07801_ (.Y(_02100_),
    .A(_02099_),
    .B(_02063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07802_ (.Y(_02101_),
    .B1(\acc_sub.exp_mant_logic0.b[2] ),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[5] ),
    .A1(net1779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07803_ (.Y(_01415_),
    .A(_02100_),
    .B(_02101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07804_ (.Y(_02102_),
    .A(_01989_),
    .B(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07805_ (.Y(_02103_),
    .A(net1650),
    .B(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07806_ (.Y(_02104_),
    .A(_02102_),
    .B(_02103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07807_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc_sub.exp_mant_logic0.b[3] ),
    .A2(net1646),
    .Y(_02105_),
    .B1(_02104_));
 sg13g2_a22oi_1 _07808_ (.Y(_02106_),
    .B1(\acc_sub.exp_mant_logic0.b[4] ),
    .B2(net1649),
    .A2(\acc_sub.exp_mant_logic0.b[2] ),
    .A1(net1651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07809_ (.Y(_02107_),
    .B1(net1794),
    .B2(_01975_),
    .A2(net1685),
    .A1(\acc_sub.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07810_ (.B(_02106_),
    .C(_02107_),
    .A(_02105_),
    .Y(_02108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07811_ (.Y(_02109_),
    .A(_02108_),
    .B(net1640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07812_ (.Y(_02110_),
    .B1(\acc_sub.exp_mant_logic0.b[1] ),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[4] ),
    .A1(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07813_ (.Y(_01414_),
    .A(_02109_),
    .B(_02110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07814_ (.Y(_02111_),
    .A(_02006_),
    .B(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07815_ (.Y(_02112_),
    .A(_01989_),
    .B(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07816_ (.Y(_02113_),
    .A(_01975_),
    .B(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07817_ (.B(_02112_),
    .C(_02113_),
    .A(_02111_),
    .Y(_02114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07818_ (.Y(_02115_),
    .A(net1649),
    .B(\acc_sub.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07819_ (.Y(_02116_),
    .A(net1646),
    .B(\acc_sub.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07820_ (.Y(_02117_),
    .A(net1650),
    .B(\acc_sub.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07821_ (.B(_02116_),
    .C(_02117_),
    .A(_02115_),
    .Y(_02118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07822_ (.A(_02114_),
    .B(_02118_),
    .Y(_02119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07823_ (.Y(_02120_),
    .B1(\acc_sub.exp_mant_logic0.b[1] ),
    .B2(net1651),
    .A2(net1685),
    .A1(\acc_sub.exp_mant_logic0.b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07824_ (.Y(_02121_),
    .A(_02119_),
    .B(_02120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07825_ (.Y(_02122_),
    .A(_02121_),
    .B(net1640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07826_ (.Y(_02123_),
    .B1(\acc_sub.exp_mant_logic0.b[0] ),
    .B2(net1669),
    .A2(\acc_sub.op_sign_logic0.mantisa_b[3] ),
    .A1(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07827_ (.Y(_01413_),
    .A(_02122_),
    .B(_02123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07828_ (.A(_02073_),
    .B(_01977_),
    .Y(_02124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07829_ (.A(_02091_),
    .B(_02015_),
    .Y(_02125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07830_ (.Y(_02126_),
    .A(_02006_),
    .B(\acc_sub.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07831_ (.Y(_02127_),
    .A(_02018_),
    .B(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07832_ (.Y(_02128_),
    .A(_02126_),
    .B(_02127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07833_ (.A(_02124_),
    .B(_02125_),
    .C(_02128_),
    .Y(_02129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07834_ (.VDD(VPWR),
    .Y(_02130_),
    .A(\acc_sub.exp_mant_logic0.b[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _07835_ (.Y(_02131_),
    .A(_01949_),
    .B(\acc_sub.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07836_ (.B1(_02131_),
    .VDD(VPWR),
    .Y(_02132_),
    .VSS(VGND),
    .A1(_02130_),
    .A2(_01979_));
 sg13g2_nand2_1 _07837_ (.Y(_02133_),
    .A(_01959_),
    .B(\acc_sub.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07838_ (.B1(_02133_),
    .VDD(VPWR),
    .Y(_02134_),
    .VSS(VGND),
    .A1(_02089_),
    .A2(_02024_));
 sg13g2_nor2_1 _07839_ (.A(_02132_),
    .B(_02134_),
    .Y(_02135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07840_ (.Y(_02136_),
    .A(_02129_),
    .B(_02135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07841_ (.Y(_02137_),
    .A(_02136_),
    .B(net1640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07842_ (.Y(_02138_),
    .A(net1779),
    .B(\acc_sub.op_sign_logic0.mantisa_b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07843_ (.Y(_01412_),
    .A(_02137_),
    .B(_02138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07844_ (.Y(_02139_),
    .A(_01959_),
    .B(\acc_sub.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07845_ (.B1(_02139_),
    .VDD(VPWR),
    .Y(_02140_),
    .VSS(VGND),
    .A1(_02073_),
    .A2(_02015_));
 sg13g2_nor2_1 _07846_ (.A(_02089_),
    .B(_01977_),
    .Y(_02141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07847_ (.Y(_02142_),
    .A(_02018_),
    .B(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07848_ (.Y(_02143_),
    .A(_02006_),
    .B(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07849_ (.Y(_02144_),
    .A(_02142_),
    .B(_02143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07850_ (.A(_02141_),
    .B(_02144_),
    .Y(_02145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07851_ (.Y(_02146_),
    .B1(\acc_sub.exp_mant_logic0.b[0] ),
    .B2(_01949_),
    .A2(\acc_sub.exp_mant_logic0.b[2] ),
    .A1(net1650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _07852_ (.B(_02145_),
    .C(_02146_),
    .Y(_02147_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_02140_));
 sg13g2_nand2_1 _07853_ (.Y(_02148_),
    .A(_02147_),
    .B(net1640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07854_ (.Y(_02149_),
    .A(net1779),
    .B(\acc_sub.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07855_ (.Y(_01411_),
    .A(_02148_),
    .B(_02149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07856_ (.Y(_02150_),
    .A(_02006_),
    .B(\acc_sub.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07857_ (.Y(_02151_),
    .A(_02018_),
    .B(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07858_ (.Y(_02152_),
    .A(_02150_),
    .B(_02151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07859_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc_sub.exp_mant_logic0.b[2] ),
    .A2(_01975_),
    .Y(_02153_),
    .B1(_02152_));
 sg13g2_nor2_1 _07860_ (.A(_02089_),
    .B(_02015_),
    .Y(_02154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07861_ (.A(_02130_),
    .B(_02048_),
    .Y(_02155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07862_ (.VDD(VPWR),
    .Y(_02156_),
    .A(\acc_sub.exp_mant_logic0.b[1] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07863_ (.A(_02156_),
    .B(_02024_),
    .Y(_02157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _07864_ (.A(_02154_),
    .B(_02155_),
    .C(_02157_),
    .Y(_02158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07865_ (.Y(_02159_),
    .A(_02153_),
    .B(_02158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07866_ (.Y(_02160_),
    .A(_02159_),
    .B(_02063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07867_ (.B1(_02160_),
    .VDD(VPWR),
    .Y(_01410_),
    .VSS(VGND),
    .A1(\acc_sub.reg1en.q[0] ),
    .A2(_01545_));
 sg13g2_nand2_1 _07868_ (.Y(_02161_),
    .A(net1885),
    .B(\acc_sub.x2[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07869_ (.B1(_02161_),
    .VDD(VPWR),
    .Y(_01409_),
    .VSS(VGND),
    .A1(net1885),
    .A2(_01776_));
 sg13g2_nand2_1 _07870_ (.Y(_02162_),
    .A(net1888),
    .B(\acc_sub.x2[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07871_ (.B1(_02162_),
    .VDD(VPWR),
    .Y(_01408_),
    .VSS(VGND),
    .A1(net1887),
    .A2(_01789_));
 sg13g2_nand2_1 _07872_ (.Y(_02163_),
    .A(net1888),
    .B(\acc_sub.x2[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07873_ (.B1(_02163_),
    .VDD(VPWR),
    .Y(_01407_),
    .VSS(VGND),
    .A1(net1889),
    .A2(_01784_));
 sg13g2_nand2_1 _07874_ (.Y(_02164_),
    .A(net1888),
    .B(\acc_sub.x2[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07875_ (.B1(_02164_),
    .VDD(VPWR),
    .Y(_01406_),
    .VSS(VGND),
    .A1(net1887),
    .A2(_01795_));
 sg13g2_nand2_1 _07876_ (.Y(_02165_),
    .A(net1888),
    .B(\acc_sub.x2[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07877_ (.B1(_02165_),
    .VDD(VPWR),
    .Y(_01405_),
    .VSS(VGND),
    .A1(net1888),
    .A2(_01799_));
 sg13g2_nand2_1 _07878_ (.Y(_02166_),
    .A(net1886),
    .B(\acc_sub.x2[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07879_ (.B1(_02166_),
    .VDD(VPWR),
    .Y(_01404_),
    .VSS(VGND),
    .A1(net1885),
    .A2(_01804_));
 sg13g2_nand2_1 _07880_ (.Y(_02167_),
    .A(net1885),
    .B(\acc_sub.x2[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07881_ (.B1(_02167_),
    .VDD(VPWR),
    .Y(_01403_),
    .VSS(VGND),
    .A1(net1895),
    .A2(_01808_));
 sg13g2_nand2_1 _07882_ (.Y(_02168_),
    .A(net1887),
    .B(\acc_sub.x2[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07883_ (.B1(_02168_),
    .VDD(VPWR),
    .Y(_01402_),
    .VSS(VGND),
    .A1(net1895),
    .A2(_01825_));
 sg13g2_nand2_1 _07884_ (.Y(_02169_),
    .A(net1888),
    .B(\acc_sub.x2[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07885_ (.B1(_02169_),
    .VDD(VPWR),
    .Y(_01401_),
    .VSS(VGND),
    .A1(net1895),
    .A2(_01813_));
 sg13g2_nand2_1 _07886_ (.Y(_02170_),
    .A(net1892),
    .B(\acc_sub.x2[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07887_ (.B1(_02170_),
    .VDD(VPWR),
    .Y(_01400_),
    .VSS(VGND),
    .A1(net1892),
    .A2(_02096_));
 sg13g2_nand2_1 _07888_ (.Y(_02171_),
    .A(net1891),
    .B(\acc_sub.x2[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07889_ (.B1(_02171_),
    .VDD(VPWR),
    .Y(_01399_),
    .VSS(VGND),
    .A1(net1891),
    .A2(_02091_));
 sg13g2_nand2_1 _07890_ (.Y(_02172_),
    .A(net1892),
    .B(\acc_sub.x2[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07891_ (.B1(_02172_),
    .VDD(VPWR),
    .Y(_01398_),
    .VSS(VGND),
    .A1(net1892),
    .A2(_02073_));
 sg13g2_nand2_1 _07892_ (.Y(_02173_),
    .A(net1892),
    .B(\acc_sub.x2[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07893_ (.B1(_02173_),
    .VDD(VPWR),
    .Y(_01397_),
    .VSS(VGND),
    .A1(net1892),
    .A2(_02089_));
 sg13g2_nand2_1 _07894_ (.Y(_02174_),
    .A(net1891),
    .B(\acc_sub.x2[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07895_ (.B1(_02174_),
    .VDD(VPWR),
    .Y(_01396_),
    .VSS(VGND),
    .A1(net1891),
    .A2(_02087_));
 sg13g2_nand2_1 _07896_ (.Y(_02175_),
    .A(net1891),
    .B(\acc_sub.x2[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07897_ (.B1(_02175_),
    .VDD(VPWR),
    .Y(_01395_),
    .VSS(VGND),
    .A1(net1891),
    .A2(_02156_));
 sg13g2_nand2_1 _07898_ (.Y(_02176_),
    .A(net1892),
    .B(\acc_sub.x2[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07899_ (.B1(_02176_),
    .VDD(VPWR),
    .Y(_01394_),
    .VSS(VGND),
    .A1(net1892),
    .A2(_02130_));
 sg13g2_mux2_1 _07900_ (.A0(\fp16_sum_pipe.op_sign_logic0.s_a ),
    .A1(\fp16_sum_pipe.exp_mant_logic0.a[15] ),
    .S(\fp16_sum_pipe.reg1en.q[0] ),
    .X(_01393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07901_ (.VDD(VPWR),
    .Y(_02177_),
    .A(\fp16_sum_pipe.op_sign_logic0.s_b ),
    .VSS(VGND));
 sg13g2_nand2_1 _07902_ (.Y(_02178_),
    .A(net1843),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07903_ (.B1(_02178_),
    .VDD(VPWR),
    .Y(_01392_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.reg1en.q[0] ),
    .A2(_02177_));
 sg13g2_inv_2 _07904_ (.Y(_02179_),
    .A(\fp16_sum_pipe.reg1en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout50 (.A(net51),
    .X(net50),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1788 (.A(\acc_sub.add_renorm0.mantisa[11] ),
    .X(net1788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07907_ (.VDD(VPWR),
    .Y(_02182_),
    .A(\fp16_sum_pipe.seg_reg0.q[29] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07908_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[14] ),
    .B(_02179_),
    .Y(_02183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _07909_ (.Y(_02184_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[14] ),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07910_ (.VDD(VPWR),
    .Y(_02185_),
    .A(_02184_),
    .VSS(VGND));
 sg13g2_inv_2 _07911_ (.Y(_02186_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07912_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[13] ),
    .B(_02186_),
    .Y(_02187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07913_ (.VDD(VPWR),
    .Y(_02188_),
    .A(_02187_),
    .VSS(VGND));
 sg13g2_nand2_1 _07914_ (.Y(_02189_),
    .A(_02186_),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07915_ (.Y(_02190_),
    .A(_02188_),
    .B(_02189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07916_ (.A(_02185_),
    .B(_02190_),
    .Y(_02191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07917_ (.VDD(VPWR),
    .Y(_02192_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[11] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07918_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[11] ),
    .B(_02192_),
    .Y(_02193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07919_ (.Y(_02194_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07920_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[11] ),
    .B(_02194_),
    .Y(_02195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07921_ (.A(_02193_),
    .B(_02195_),
    .Y(_02196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07922_ (.Y(_02197_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07923_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[12] ),
    .B(_02197_),
    .Y(_02198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _07924_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[12] ),
    .Y(_02199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07925_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[12] ),
    .B(_02199_),
    .Y(_02200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07926_ (.A(_02198_),
    .B(_02200_),
    .Y(_02201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _07927_ (.X(_02202_),
    .A(_02191_),
    .B(_02196_),
    .C(_02201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07928_ (.VDD(VPWR),
    .Y(_02203_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07929_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[10] ),
    .B(_02203_),
    .Y(_02204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07930_ (.Y(_02205_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07931_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[10] ),
    .B(_02205_),
    .Y(_02206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07932_ (.A(_02204_),
    .B(_02206_),
    .Y(_02207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07933_ (.VDD(VPWR),
    .Y(_02208_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[9] ),
    .VSS(VGND));
 sg13g2_nor2_1 _07934_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[9] ),
    .B(_02208_),
    .Y(_02209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07935_ (.Y(_02210_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07936_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[9] ),
    .B(_02210_),
    .Y(_02211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07937_ (.A(_02209_),
    .B(_02211_),
    .Y(_02212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07938_ (.Y(_02213_),
    .A(_02207_),
    .B(_02212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _07939_ (.B(\fp16_sum_pipe.exp_mant_logic0.b[8] ),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[8] ),
    .X(_02214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07940_ (.VDD(VPWR),
    .Y(_02215_),
    .A(_02214_),
    .VSS(VGND));
 sg13g2_inv_2 _07941_ (.Y(_02216_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07942_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[7] ),
    .B(_02216_),
    .Y(_02217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07943_ (.Y(_02218_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07944_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[7] ),
    .B(_02218_),
    .Y(_02219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07945_ (.A(_02217_),
    .B(_02219_),
    .Y(_02220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07946_ (.Y(_02221_),
    .A(_02215_),
    .B(_02220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07947_ (.A(_02213_),
    .B(_02221_),
    .Y(_02222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _07948_ (.Y(_02223_),
    .A(_02202_),
    .B(_02222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout121 (.A(net122),
    .X(net121),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07950_ (.Y(_02225_),
    .A(_02223_),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07951_ (.Y(_01391_),
    .B1(_02183_),
    .B2(_02225_),
    .A2(_02182_),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07952_ (.VDD(VPWR),
    .Y(_02226_),
    .A(\fp16_sum_pipe.seg_reg0.q[28] ),
    .VSS(VGND));
 sg13g2_inv_2 _07953_ (.Y(_02227_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _07954_ (.Y(_02228_),
    .A(_02227_),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07955_ (.B1(_02228_),
    .VDD(VPWR),
    .Y(_02229_),
    .VSS(VGND),
    .A1(_02217_),
    .A2(_02214_));
 sg13g2_inv_1 _07956_ (.VDD(VPWR),
    .Y(_02230_),
    .A(_02211_),
    .VSS(VGND));
 sg13g2_a21oi_1 _07957_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02229_),
    .A2(_02230_),
    .Y(_02231_),
    .B1(_02209_));
 sg13g2_inv_1 _07958_ (.VDD(VPWR),
    .Y(_02232_),
    .A(_02204_),
    .VSS(VGND));
 sg13g2_o21ai_1 _07959_ (.B1(_02232_),
    .VDD(VPWR),
    .Y(_02233_),
    .VSS(VGND),
    .A1(_02206_),
    .A2(_02231_));
 sg13g2_nand2_1 _07960_ (.Y(_02234_),
    .A(_02233_),
    .B(_02202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _07961_ (.VDD(VPWR),
    .Y(_02235_),
    .A(_02193_),
    .VSS(VGND));
 sg13g2_inv_1 _07962_ (.VDD(VPWR),
    .Y(_02236_),
    .A(_02198_),
    .VSS(VGND));
 sg13g2_o21ai_1 _07963_ (.B1(_02236_),
    .VDD(VPWR),
    .Y(_02237_),
    .VSS(VGND),
    .A1(_02200_),
    .A2(_02235_));
 sg13g2_inv_2 _07964_ (.Y(_02238_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _07965_ (.A(\fp16_sum_pipe.exp_mant_logic0.b[14] ),
    .B(_02238_),
    .Y(_02239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _07966_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02191_),
    .C1(_02239_),
    .B1(_02237_),
    .A1(_02187_),
    .Y(_02240_),
    .A2(_02184_));
 sg13g2_nand2_2 _07967_ (.Y(_02241_),
    .A(_02234_),
    .B(_02240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _07968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02241_),
    .A2(_02186_),
    .Y(_02242_),
    .B1(_02179_));
 sg13g2_o21ai_1 _07969_ (.B1(_02242_),
    .VDD(VPWR),
    .Y(_02243_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.exp_mant_logic0.b[13] ),
    .A2(_02241_));
 sg13g2_o21ai_1 _07970_ (.B1(_02243_),
    .VDD(VPWR),
    .Y(_01390_),
    .VSS(VGND),
    .A1(net1843),
    .A2(_02226_));
 sg13g2_nand2_2 _07971_ (.Y(_02244_),
    .A(_02241_),
    .B(_02223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _07972_ (.A(_02244_),
    .Y(_02245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07973_ (.A(_02179_),
    .B(_02245_),
    .Y(_02246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _07975_ (.A(_02246_),
    .Y(_02248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1703 (.A(_04029_),
    .X(net1703),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _07977_ (.A(_02179_),
    .B(_02244_),
    .Y(_02250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _07980_ (.Y(_02253_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[12] ),
    .B2(_02250_),
    .A2(\fp16_sum_pipe.seg_reg0.q[27] ),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07981_ (.B1(_02253_),
    .VDD(VPWR),
    .Y(_01389_),
    .VSS(VGND),
    .A1(_02199_),
    .A2(_02248_));
 sg13g2_a22oi_1 _07982_ (.Y(_02254_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[11] ),
    .B2(_02250_),
    .A2(\fp16_sum_pipe.seg_reg0.q[26] ),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07983_ (.B1(_02254_),
    .VDD(VPWR),
    .Y(_01388_),
    .VSS(VGND),
    .A1(_02194_),
    .A2(_02248_));
 sg13g2_a22oi_1 _07984_ (.Y(_02255_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[10] ),
    .B2(_02250_),
    .A2(\fp16_sum_pipe.seg_reg0.q[25] ),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07985_ (.B1(_02255_),
    .VDD(VPWR),
    .Y(_01387_),
    .VSS(VGND),
    .A1(_02205_),
    .A2(_02248_));
 sg13g2_a22oi_1 _07986_ (.Y(_02256_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[9] ),
    .B2(_02250_),
    .A2(\fp16_sum_pipe.seg_reg0.q[24] ),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07987_ (.B1(_02256_),
    .VDD(VPWR),
    .Y(_01386_),
    .VSS(VGND),
    .A1(_02210_),
    .A2(_02248_));
 sg13g2_a22oi_1 _07988_ (.Y(_02257_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[8] ),
    .B2(_02250_),
    .A2(\fp16_sum_pipe.seg_reg0.q[23] ),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07989_ (.B1(_02257_),
    .VDD(VPWR),
    .Y(_01385_),
    .VSS(VGND),
    .A1(_02227_),
    .A2(_02248_));
 sg13g2_a22oi_1 _07990_ (.Y(_02258_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[7] ),
    .B2(_02250_),
    .A2(\fp16_sum_pipe.seg_reg0.q[22] ),
    .A1(net1775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _07991_ (.B1(_02258_),
    .VDD(VPWR),
    .Y(_01384_),
    .VSS(VGND),
    .A1(_02216_),
    .A2(_02248_));
 sg13g2_inv_1 _07992_ (.VDD(VPWR),
    .Y(_02259_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[10] ),
    .VSS(VGND));
 sg13g2_inv_2 _07993_ (.Y(_02260_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _07994_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .Y(_02261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07995_ (.Y(_02262_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _07996_ (.B(_02261_),
    .C(_02262_),
    .A(_02260_),
    .Y(_02263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _07997_ (.Y(_02264_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _07998_ (.B(_02208_),
    .C(_02264_),
    .A(_02203_),
    .Y(_02265_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02218_));
 sg13g2_nand4_1 _07999_ (.B(_02186_),
    .C(_02197_),
    .A(_02238_),
    .Y(_02266_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02192_));
 sg13g2_inv_2 _08000_ (.Y(_02267_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08001_ (.Y(_02268_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _08002_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[2] ),
    .Y(_02269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08003_ (.Y(_02270_),
    .A(\fp16_sum_pipe.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08004_ (.B(_02268_),
    .C(_02269_),
    .A(_02267_),
    .Y(_02271_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02270_));
 sg13g2_nor4_2 _08005_ (.A(_02263_),
    .B(_02265_),
    .C(_02266_),
    .Y(_02272_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_02271_));
 sg13g2_inv_4 _08006_ (.A(_02272_),
    .Y(_02273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08007_ (.B(net1843),
    .C(_02273_),
    .A(_02241_),
    .Y(_02274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08008_ (.B1(_02274_),
    .VDD(VPWR),
    .Y(_01383_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.reg1en.q[0] ),
    .A2(_02259_));
 sg13g2_inv_2 _08009_ (.Y(_02275_),
    .A(_02223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1719 (.A(_07076_),
    .X(net1719),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08011_ (.Y(_02277_),
    .A(_02264_),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08012_ (.B1(_02277_),
    .VDD(VPWR),
    .Y(_02278_),
    .VSS(VGND),
    .A1(_02219_),
    .A2(_02214_));
 sg13g2_inv_1 _08013_ (.VDD(VPWR),
    .Y(_02279_),
    .A(_02278_),
    .VSS(VGND));
 sg13g2_nor2_1 _08014_ (.A(_02213_),
    .B(_02279_),
    .Y(_02280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08015_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02232_),
    .A2(_02211_),
    .Y(_02281_),
    .B1(_02206_));
 sg13g2_nor2b_1 _08016_ (.A(_02280_),
    .B_N(_02281_),
    .Y(_02282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08017_ (.VDD(VPWR),
    .Y(_02283_),
    .A(_02282_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08018_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02283_),
    .A2(_02235_),
    .Y(_02284_),
    .B1(_02195_));
 sg13g2_inv_1 _08019_ (.VDD(VPWR),
    .Y(_02285_),
    .A(_02284_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08020_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02285_),
    .A2(_02236_),
    .Y(_02286_),
    .B1(_02200_));
 sg13g2_a21o_1 _08021_ (.A2(_02189_),
    .A1(_02286_),
    .B1(_02187_),
    .X(_02287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08022_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02233_),
    .A2(_02196_),
    .Y(_02288_),
    .B1(_02193_));
 sg13g2_o21ai_1 _08023_ (.B1(_02236_),
    .VDD(VPWR),
    .Y(_02289_),
    .VSS(VGND),
    .A1(_02200_),
    .A2(_02288_));
 sg13g2_nand2_1 _08024_ (.Y(_02290_),
    .A(_02289_),
    .B(_02189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08025_ (.Y(_02291_),
    .B1(_02188_),
    .B2(_02290_),
    .A2(\fp16_sum_pipe.exp_mant_logic0.b[14] ),
    .A1(_02238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08026_ (.Y(_02292_),
    .A(_02291_),
    .B(_02223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08027_ (.B1(_02292_),
    .VDD(VPWR),
    .Y(_02293_),
    .VSS(VGND),
    .A1(_02245_),
    .A2(_02287_));
 sg13g2_nand2_1 _08028_ (.Y(_02294_),
    .A(_02293_),
    .B(_02185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08029_ (.A(_02233_),
    .B(net1692),
    .Y(_02295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1692),
    .A2(_02282_),
    .Y(_02296_),
    .B1(_02295_));
 sg13g2_xor2_1 _08031_ (.B(_02296_),
    .A(_02196_),
    .X(_02297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08032_ (.Y(_02298_),
    .A(net1692),
    .B(_02285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08033_ (.B1(_02298_),
    .VDD(VPWR),
    .Y(_02299_),
    .VSS(VGND),
    .A1(_02288_),
    .A2(net1692));
 sg13g2_xor2_1 _08034_ (.B(_02299_),
    .A(_02201_),
    .X(_02300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08035_ (.A(_02286_),
    .B(_02245_),
    .Y(_02301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08036_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02289_),
    .A2(_02245_),
    .Y(_02302_),
    .B1(_02301_));
 sg13g2_xor2_1 _08037_ (.B(_02302_),
    .A(_02190_),
    .X(_02303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08038_ (.A(_02297_),
    .B(_02300_),
    .C(_02303_),
    .Y(_02304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08039_ (.Y(_02305_),
    .A(_02294_),
    .B(_02304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1818 (.A(net1816),
    .X(net1818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08041_ (.Y(_02307_),
    .A(_02305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08042_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02279_),
    .A2(_02230_),
    .Y(_02308_),
    .B1(_02209_));
 sg13g2_nor2_1 _08043_ (.A(_02308_),
    .B(_02245_),
    .Y(_02309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08044_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02231_),
    .A2(_02245_),
    .Y(_02310_),
    .B1(_02309_));
 sg13g2_xnor2_1 _08045_ (.Y(_02311_),
    .A(_02207_),
    .B(_02310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08046_ (.Y(_02312_),
    .A(net1692),
    .B(_02279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08047_ (.B1(_02312_),
    .VDD(VPWR),
    .Y(_02313_),
    .VSS(VGND),
    .A1(_02229_),
    .A2(net1692));
 sg13g2_xor2_1 _08048_ (.B(_02313_),
    .A(_02212_),
    .X(_02314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08049_ (.Y(_02315_),
    .A(_02311_),
    .B(_02314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08050_ (.Y(_02316_),
    .B(net1692),
    .A_N(_02219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08051_ (.B1(_02316_),
    .VDD(VPWR),
    .Y(_02317_),
    .VSS(VGND),
    .A1(_02217_),
    .A2(net1692));
 sg13g2_xnor2_1 _08052_ (.Y(_02318_),
    .A(_02214_),
    .B(_02317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08053_ (.VDD(VPWR),
    .Y(_02319_),
    .A(_02220_),
    .VSS(VGND));
 sg13g2_nand2b_1 _08054_ (.Y(_02320_),
    .B(_02319_),
    .A_N(_02318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08055_ (.A(_02315_),
    .B(_02320_),
    .Y(_02321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08056_ (.Y(_02322_),
    .A(_02307_),
    .B(_02321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_74_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_74_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08058_ (.VDD(VPWR),
    .Y(_02324_),
    .A(net1652),
    .VSS(VGND));
 sg13g2_a22oi_1 _08059_ (.Y(_02325_),
    .B1(_02273_),
    .B2(_02324_),
    .A2(net1691),
    .A1(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08060_ (.VDD(VPWR),
    .Y(_02326_),
    .A(_02314_),
    .VSS(VGND));
 sg13g2_nand2_2 _08061_ (.Y(_02327_),
    .A(_02311_),
    .B(_02326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08062_ (.VDD(VPWR),
    .Y(_02328_),
    .A(_02327_),
    .VSS(VGND));
 sg13g2_nand2_1 _08063_ (.Y(_02329_),
    .A(_02328_),
    .B(_02221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08064_ (.B1(_02223_),
    .VDD(VPWR),
    .Y(_02330_),
    .VSS(VGND),
    .A1(_02329_),
    .A2(_02305_));
 sg13g2_nor3_1 _08065_ (.A(_02221_),
    .B(_02326_),
    .C(_02311_),
    .Y(_02331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08066_ (.A(_02305_),
    .B_N(_02331_),
    .Y(_02332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1664 (.A(_03681_),
    .X(net1664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08068_ (.VDD(VPWR),
    .Y(_02334_),
    .A(_02332_),
    .VSS(VGND));
 sg13g2_nand2_1 _08069_ (.Y(_02335_),
    .A(_02334_),
    .B(net1652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08070_ (.Y(_02336_),
    .A(_02220_),
    .B(_02214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08071_ (.A(_02336_),
    .B(_02315_),
    .Y(_02337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08072_ (.A(_02305_),
    .B_N(_02337_),
    .Y(_02338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_57_clk (.A(clknet_5_25__leaf_clk),
    .X(clknet_leaf_57_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08074_ (.Y(_02340_),
    .A(_02338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08075_ (.Y(_02341_),
    .A(_02318_),
    .B(_02319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08076_ (.A(_02341_),
    .B(_02315_),
    .Y(_02342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08077_ (.A(_02305_),
    .B_N(_02342_),
    .Y(_02343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1663 (.A(_05106_),
    .X(net1663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08079_ (.Y(_02345_),
    .A(_02343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08080_ (.A(_02221_),
    .B(_02327_),
    .Y(_02346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08081_ (.A(_02305_),
    .B_N(_02346_),
    .Y(_02347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_59_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_59_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08083_ (.Y(_02349_),
    .A(_02347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08084_ (.B(_02345_),
    .C(_02349_),
    .A(_02340_),
    .Y(_02350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08085_ (.A(_02330_),
    .B(_02335_),
    .C(_02350_),
    .Y(_02351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08086_ (.A(_02248_),
    .B(_02351_),
    .Y(_02352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_97_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_97_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08088_ (.Y(_02354_),
    .B(net1639),
    .A_N(_02325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08089_ (.Y(_02355_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[9] ),
    .A1(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08090_ (.Y(_01382_),
    .A(_02354_),
    .B(_02355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08091_ (.Y(_02356_),
    .A(net1645),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_56_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_56_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08093_ (.Y(_02358_),
    .A(net1659),
    .B(_02273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08094_ (.Y(_02359_),
    .A(net1691),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08095_ (.B(_02358_),
    .C(_02359_),
    .A(_02356_),
    .Y(_02360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08096_ (.Y(_02361_),
    .A(net1639),
    .B(_02360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08097_ (.Y(_02362_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[8] ),
    .A1(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08098_ (.Y(_01381_),
    .A(_02361_),
    .B(_02362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08099_ (.Y(_02363_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .B2(net1659),
    .A2(net1691),
    .A1(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08100_ (.Y(_02364_),
    .A(net1645),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08101_ (.Y(_02365_),
    .A(_02343_),
    .B(_02273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08102_ (.B(_02364_),
    .C(_02365_),
    .A(_02363_),
    .Y(_02366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08103_ (.Y(_02367_),
    .A(net1639),
    .B(_02366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout49 (.A(net72),
    .X(net49),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08105_ (.Y(_02369_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[7] ),
    .A1(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08106_ (.Y(_01380_),
    .A(_02367_),
    .B(_02369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08107_ (.Y(_02370_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .B2(net1645),
    .A2(_02343_),
    .A1(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08108_ (.Y(_02371_),
    .A(net1658),
    .B(_02273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08109_ (.Y(_02372_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .B2(net1659),
    .A2(net1691),
    .A1(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08110_ (.B(_02371_),
    .C(_02372_),
    .A(_02370_),
    .Y(_02373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08111_ (.Y(_02374_),
    .A(net1639),
    .B(_02373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08112_ (.Y(_02375_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[6] ),
    .A1(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08113_ (.Y(_01379_),
    .A(_02374_),
    .B(_02375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08114_ (.A(_02268_),
    .B(net1652),
    .Y(_02376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08115_ (.A(_02327_),
    .B(_02320_),
    .Y(_02377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08116_ (.A(_02305_),
    .B_N(_02377_),
    .Y(_02378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_61_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_61_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08118_ (.Y(_02380_),
    .A(net1657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08119_ (.A(_02272_),
    .B(_02380_),
    .Y(_02381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_90_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_90_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08121_ (.A(_02260_),
    .B(net1648),
    .Y(_02383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08122_ (.A(_02376_),
    .B(_02381_),
    .C(_02383_),
    .Y(_02384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08123_ (.A(_02269_),
    .B(_02223_),
    .Y(_02385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08124_ (.A(_02261_),
    .B(_02340_),
    .Y(_02386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08125_ (.A(_02267_),
    .B(_02349_),
    .Y(_02387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08126_ (.A(_02385_),
    .B(_02386_),
    .C(_02387_),
    .Y(_02388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08127_ (.Y(_02389_),
    .A(_02384_),
    .B(_02388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08128_ (.Y(_02390_),
    .A(_02352_),
    .B(_02389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08129_ (.Y(_02391_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[2] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[5] ),
    .A1(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08130_ (.Y(_01378_),
    .A(_02390_),
    .B(_02391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08131_ (.A(_02269_),
    .B(net1652),
    .Y(_02392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08132_ (.A(_02261_),
    .B(net1648),
    .Y(_02393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08133_ (.A(_02267_),
    .B(_02380_),
    .Y(_02394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08134_ (.A(_02392_),
    .B(_02393_),
    .C(_02394_),
    .Y(_02395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _08135_ (.B(_02307_),
    .C(_02328_),
    .Y(_02396_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_02336_));
 sg13g2_buf_2 place1657 (.A(_02378_),
    .X(net1657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08137_ (.A(_02272_),
    .B(_02396_),
    .Y(_02398_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08138_ (.Y(_02399_),
    .A(net1691),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08139_ (.A(_02398_),
    .B_N(_02399_),
    .Y(_02400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08140_ (.Y(_02401_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .B2(net1658),
    .A2(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .A1(net1659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08141_ (.B(_02400_),
    .C(_02401_),
    .A(_02395_),
    .Y(_02402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08142_ (.Y(_02403_),
    .A(_02402_),
    .B(_02352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08143_ (.Y(_02404_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[1] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[4] ),
    .A1(net1774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08144_ (.Y(_01377_),
    .A(_02403_),
    .B(_02404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08145_ (.Y(_02405_),
    .A(_02378_),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08146_ (.B1(_02405_),
    .VDD(VPWR),
    .Y(_02406_),
    .VSS(VGND),
    .A1(_02262_),
    .A2(net1652));
 sg13g2_nor2_1 _08147_ (.A(_02341_),
    .B(_02327_),
    .Y(_02407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08148_ (.A(_02305_),
    .B_N(_02407_),
    .Y(_02408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1661 (.A(_05146_),
    .X(net1661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08150_ (.Y(_02410_),
    .A(_02408_),
    .B(_02273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08151_ (.B1(_02410_),
    .VDD(VPWR),
    .Y(_02411_),
    .VSS(VGND),
    .A1(_02268_),
    .A2(net1648));
 sg13g2_nor2_1 _08152_ (.A(_02406_),
    .B(_02411_),
    .Y(_02412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08153_ (.Y(_02413_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .B2(net1658),
    .A2(net1691),
    .A1(\fp16_sum_pipe.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08154_ (.A(_02267_),
    .B(_02396_),
    .Y(_02414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08155_ (.Y(_02415_),
    .A(net1659),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08156_ (.A(_02414_),
    .B_N(_02415_),
    .Y(_02416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08157_ (.B(_02413_),
    .C(_02416_),
    .A(_02412_),
    .Y(_02417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08158_ (.Y(_02418_),
    .A(_02417_),
    .B(net1639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08159_ (.Y(_02419_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[0] ),
    .B2(net1684),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_a[3] ),
    .A1(net1776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08160_ (.Y(_01376_),
    .A(_02418_),
    .B(_02419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08161_ (.Y(_02420_),
    .A(net1659),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08162_ (.B1(_02420_),
    .VDD(VPWR),
    .Y(_02421_),
    .VSS(VGND),
    .A1(_02270_),
    .A2(net1652));
 sg13g2_nand2_1 _08163_ (.Y(_02422_),
    .A(net1658),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08164_ (.B1(_02422_),
    .VDD(VPWR),
    .Y(_02423_),
    .VSS(VGND),
    .A1(_02269_),
    .A2(net1648));
 sg13g2_nor2_1 _08165_ (.A(_02421_),
    .B(_02423_),
    .Y(_02424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08166_ (.Y(_02425_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .B2(_02408_),
    .A2(_02273_),
    .A1(_02332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08167_ (.A(_02336_),
    .B(_02327_),
    .Y(_02426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08168_ (.Y(_02427_),
    .A(_02307_),
    .B(_02426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08169_ (.A(_02260_),
    .B(_02427_),
    .Y(_02428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08170_ (.Y(_02429_),
    .A(_02378_),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08171_ (.A(_02428_),
    .B_N(_02429_),
    .Y(_02430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08172_ (.B(_02425_),
    .C(_02430_),
    .A(_02424_),
    .Y(_02431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08173_ (.Y(_02432_),
    .A(_02431_),
    .B(net1639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08174_ (.Y(_02433_),
    .A(net1774),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08175_ (.Y(_01375_),
    .A(_02432_),
    .B(_02433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08176_ (.A(_02270_),
    .B(_02340_),
    .Y(_02434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08177_ (.A(_02269_),
    .B(_02349_),
    .Y(_02435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08178_ (.A(_02262_),
    .B(net1648),
    .Y(_02436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08179_ (.A(_02434_),
    .B(_02435_),
    .C(_02436_),
    .Y(_02437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08180_ (.Y(_02438_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .B2(_02408_),
    .A2(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .A1(_02332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08181_ (.A(_02261_),
    .B(_02427_),
    .Y(_02439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08182_ (.Y(_02440_),
    .A(_02378_),
    .B(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08183_ (.A(_02439_),
    .B_N(_02440_),
    .Y(_02441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08184_ (.B(_02438_),
    .C(_02441_),
    .A(_02437_),
    .Y(_02442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08185_ (.Y(_02443_),
    .A(_02442_),
    .B(net1639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08186_ (.Y(_02444_),
    .A(net1774),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08187_ (.Y(_01374_),
    .A(_02443_),
    .B(_02444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08188_ (.A(_02260_),
    .B(_02334_),
    .Y(_02445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08189_ (.A(_02262_),
    .B(_02349_),
    .Y(_02446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08190_ (.A(_02268_),
    .B(_02396_),
    .Y(_02447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08191_ (.A(_02445_),
    .B(_02446_),
    .C(_02447_),
    .Y(_02448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08192_ (.A(_02269_),
    .B(_02380_),
    .Y(_02449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08193_ (.VDD(VPWR),
    .Y(_02450_),
    .A(_02408_),
    .VSS(VGND));
 sg13g2_nor2_1 _08194_ (.A(_02261_),
    .B(_02450_),
    .Y(_02451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08195_ (.A(_02270_),
    .B(net1648),
    .Y(_02452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08196_ (.A(_02449_),
    .B(_02451_),
    .C(_02452_),
    .Y(_02453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08197_ (.Y(_02454_),
    .A(_02448_),
    .B(_02453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08198_ (.Y(_02455_),
    .A(net1639),
    .B(_02454_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08199_ (.Y(_02456_),
    .A(net1774),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08200_ (.Y(_01373_),
    .A(_02455_),
    .B(_02456_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08201_ (.VDD(VPWR),
    .Y(_02457_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[10] ),
    .VSS(VGND));
 sg13g2_inv_1 _08202_ (.VDD(VPWR),
    .Y(_02458_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[5] ),
    .VSS(VGND));
 sg13g2_inv_2 _08203_ (.Y(_02459_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08204_ (.Y(_02460_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08205_ (.B(_02459_),
    .C(_02460_),
    .A(_02458_),
    .Y(_02461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08206_ (.B(_02210_),
    .C(_02227_),
    .A(_02205_),
    .Y(_02462_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02216_));
 sg13g2_inv_1 _08207_ (.VDD(VPWR),
    .Y(_02463_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[14] ),
    .VSS(VGND));
 sg13g2_inv_1 _08208_ (.VDD(VPWR),
    .Y(_02464_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[13] ),
    .VSS(VGND));
 sg13g2_nand4_1 _08209_ (.B(_02464_),
    .C(_02199_),
    .A(_02463_),
    .Y(_02465_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02194_));
 sg13g2_inv_2 _08210_ (.Y(_02466_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08211_ (.Y(_02467_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08212_ (.Y(_02468_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08213_ (.Y(_02469_),
    .A(\fp16_sum_pipe.exp_mant_logic0.b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08214_ (.B(_02467_),
    .C(_02468_),
    .A(_02466_),
    .Y(_02470_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02469_));
 sg13g2_nor4_2 _08215_ (.A(_02461_),
    .B(_02462_),
    .C(_02465_),
    .Y(_02471_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_02470_));
 sg13g2_inv_4 _08216_ (.A(_02471_),
    .Y(_02472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08217_ (.B(net1843),
    .C(_02472_),
    .A(_02244_),
    .Y(_02473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08218_ (.B1(_02473_),
    .VDD(VPWR),
    .Y(_01372_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.reg1en.q[0] ),
    .A2(_02457_));
 sg13g2_a22oi_1 _08219_ (.Y(_02474_),
    .B1(_02472_),
    .B2(net1645),
    .A2(net1691),
    .A1(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08220_ (.A(_02351_),
    .B_N(_02250_),
    .Y(_02475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_98_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_98_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08222_ (.Y(_02477_),
    .B(net1638),
    .A_N(_02474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08223_ (.Y(_02478_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[9] ),
    .A1(net1777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08224_ (.Y(_01371_),
    .A(_02477_),
    .B(_02478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08225_ (.Y(_02479_),
    .A(net1645),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08226_ (.Y(_02480_),
    .A(_02338_),
    .B(_02472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08227_ (.Y(_02481_),
    .A(net1691),
    .B(net1842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08228_ (.B(_02480_),
    .C(_02481_),
    .A(_02479_),
    .Y(_02482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08229_ (.Y(_02483_),
    .A(net1638),
    .B(_02482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08230_ (.Y(_02484_),
    .B1(net1842),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[8] ),
    .A1(net1777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08231_ (.Y(_01370_),
    .A(_02483_),
    .B(_02484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08232_ (.Y(_02485_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .B2(_02338_),
    .A2(_02275_),
    .A1(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08233_ (.Y(_02486_),
    .A(net1645),
    .B(net1842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08234_ (.Y(_02487_),
    .A(_02343_),
    .B(_02472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08235_ (.B(_02486_),
    .C(_02487_),
    .A(_02485_),
    .Y(_02488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08236_ (.Y(_02489_),
    .A(net1638),
    .B(_02488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08237_ (.Y(_02490_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[7] ),
    .A1(net1778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08238_ (.Y(_01369_),
    .A(_02489_),
    .B(_02490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08239_ (.Y(_02491_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .B2(net1645),
    .A2(_02343_),
    .A1(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08240_ (.Y(_02492_),
    .A(net1658),
    .B(_02472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08241_ (.Y(_02493_),
    .B1(net1842),
    .B2(_02338_),
    .A2(_02275_),
    .A1(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08242_ (.B(_02492_),
    .C(_02493_),
    .A(_02491_),
    .Y(_02494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08243_ (.Y(_02495_),
    .A(net1638),
    .B(_02494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08244_ (.Y(_02496_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[6] ),
    .A1(net1777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08245_ (.Y(_01368_),
    .A(_02495_),
    .B(_02496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08246_ (.A(_02468_),
    .B(_02223_),
    .Y(_02497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08247_ (.A(_02466_),
    .B(_02349_),
    .Y(_02498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08248_ (.A(_02459_),
    .B(_02340_),
    .Y(_02499_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08249_ (.A(_02497_),
    .B(_02498_),
    .C(_02499_),
    .Y(_02500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08250_ (.Y(_02501_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .B2(net1645),
    .A2(_02472_),
    .A1(net1657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08251_ (.Y(_02502_),
    .A(_02343_),
    .B(net1842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08252_ (.B(_02501_),
    .C(_02502_),
    .A(_02500_),
    .Y(_02503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08253_ (.Y(_02504_),
    .A(net1638),
    .B(_02503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08254_ (.Y(_02505_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[2] ),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[5] ),
    .A1(net1777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08255_ (.Y(_01367_),
    .A(_02504_),
    .B(_02505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08256_ (.A(_02468_),
    .B(_02322_),
    .Y(_02506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08257_ (.A(_02466_),
    .B(_02380_),
    .Y(_02507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08258_ (.A(_02459_),
    .B(_02345_),
    .Y(_02508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08259_ (.A(_02506_),
    .B(_02507_),
    .C(_02508_),
    .Y(_02509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08260_ (.A(_02471_),
    .B(_02396_),
    .Y(_02510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08261_ (.Y(_02511_),
    .A(_02347_),
    .B(net1842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08262_ (.A(_02510_),
    .B_N(_02511_),
    .Y(_02512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08263_ (.Y(_02513_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .B2(_02338_),
    .A2(_02275_),
    .A1(\fp16_sum_pipe.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08264_ (.B(_02512_),
    .C(_02513_),
    .A(_02509_),
    .Y(_02514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08265_ (.Y(_02515_),
    .A(_02514_),
    .B(_02475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08266_ (.Y(_02516_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[1] ),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[4] ),
    .A1(net1778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08267_ (.Y(_01366_),
    .A(_02515_),
    .B(_02516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08268_ (.Y(_02517_),
    .A(net1657),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08269_ (.B1(_02517_),
    .VDD(VPWR),
    .Y(_02518_),
    .VSS(VGND),
    .A1(_02460_),
    .A2(_02322_));
 sg13g2_nand2_1 _08270_ (.Y(_02519_),
    .A(_02408_),
    .B(_02472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08271_ (.B1(_02519_),
    .VDD(VPWR),
    .Y(_02520_),
    .VSS(VGND),
    .A1(_02467_),
    .A2(_02345_));
 sg13g2_nor2_1 _08272_ (.A(_02518_),
    .B(_02520_),
    .Y(_02521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08273_ (.A(_02466_),
    .B(_02396_),
    .Y(_02522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08274_ (.Y(_02523_),
    .A(_02275_),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08275_ (.A(_02522_),
    .B_N(_02523_),
    .Y(_02524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08276_ (.Y(_02525_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .B2(net1658),
    .A2(\fp16_sum_pipe.exp_mant_logic0.b[2] ),
    .A1(_02338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08277_ (.B(_02524_),
    .C(_02525_),
    .A(_02521_),
    .Y(_02526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08278_ (.Y(_02527_),
    .A(_02526_),
    .B(_02475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08279_ (.Y(_02528_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[0] ),
    .B2(_02246_),
    .A2(\fp16_sum_pipe.op_sign_logic0.mantisa_b[3] ),
    .A1(net1778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08280_ (.Y(_01365_),
    .A(_02527_),
    .B(_02528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08281_ (.Y(_02529_),
    .A(_02338_),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08282_ (.B1(_02529_),
    .VDD(VPWR),
    .Y(_02530_),
    .VSS(VGND),
    .A1(_02469_),
    .A2(_02322_));
 sg13g2_nand2_1 _08283_ (.Y(_02531_),
    .A(net1658),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08284_ (.B1(_02531_),
    .VDD(VPWR),
    .Y(_02532_),
    .VSS(VGND),
    .A1(_02468_),
    .A2(_02345_));
 sg13g2_nor2_1 _08285_ (.A(_02530_),
    .B(_02532_),
    .Y(_02533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08286_ (.Y(_02534_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .B2(_02408_),
    .A2(_02472_),
    .A1(_02332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08287_ (.A(_02458_),
    .B(_02427_),
    .Y(_02535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08288_ (.Y(_02536_),
    .A(net1657),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08289_ (.A(_02535_),
    .B_N(_02536_),
    .Y(_02537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08290_ (.B(_02534_),
    .C(_02537_),
    .A(_02533_),
    .Y(_02538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08291_ (.Y(_02539_),
    .A(_02538_),
    .B(net1638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08292_ (.Y(_02540_),
    .A(net1778),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08293_ (.Y(_01364_),
    .A(_02539_),
    .B(_02540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08294_ (.A(_02469_),
    .B(_02340_),
    .Y(_02541_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08295_ (.A(_02468_),
    .B(_02349_),
    .Y(_02542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08296_ (.A(_02460_),
    .B(_02345_),
    .Y(_02543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08297_ (.A(_02541_),
    .B(_02542_),
    .C(_02543_),
    .Y(_02544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08298_ (.Y(_02545_),
    .B1(net1842),
    .B2(_02408_),
    .A2(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .A1(_02332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08299_ (.A(_02459_),
    .B(_02427_),
    .Y(_02546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08300_ (.Y(_02547_),
    .A(net1657),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08301_ (.A(_02546_),
    .B_N(_02547_),
    .Y(_02548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08302_ (.B(_02545_),
    .C(_02548_),
    .A(_02544_),
    .Y(_02549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08303_ (.Y(_02550_),
    .A(_02549_),
    .B(net1638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08304_ (.Y(_02551_),
    .A(net1774),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08305_ (.Y(_01363_),
    .A(_02550_),
    .B(_02551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08306_ (.Y(_02552_),
    .A(net1657),
    .B(\fp16_sum_pipe.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08307_ (.B1(_02552_),
    .VDD(VPWR),
    .Y(_02553_),
    .VSS(VGND),
    .A1(_02467_),
    .A2(_02427_));
 sg13g2_a22oi_1 _08308_ (.Y(_02554_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .B2(_02408_),
    .A2(net1842),
    .A1(_02332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08309_ (.Y(_02555_),
    .B1(\fp16_sum_pipe.exp_mant_logic0.b[1] ),
    .B2(net1658),
    .A2(\fp16_sum_pipe.exp_mant_logic0.b[0] ),
    .A1(_02343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _08310_ (.B(_02554_),
    .C(_02555_),
    .Y(_02556_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_02553_));
 sg13g2_nand2_1 _08311_ (.Y(_02557_),
    .A(net1638),
    .B(_02556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08312_ (.Y(_02558_),
    .A(net1778),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08313_ (.Y(_01362_),
    .A(_02557_),
    .B(_02558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08314_ (.Y(_02559_),
    .A(\state[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08315_ (.Y(_02560_),
    .A(\state[1] ),
    .B(\state[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08316_ (.A(\state[3] ),
    .B(\state[2] ),
    .Y(_02561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08317_ (.VDD(VPWR),
    .Y(_02562_),
    .A(_02561_),
    .VSS(VGND));
 sg13g2_nor2_2 _08318_ (.A(_02560_),
    .B(_02562_),
    .Y(_02563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08319_ (.A(\state[1] ),
    .B(\state[0] ),
    .Y(_02564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08320_ (.Y(_02565_),
    .A(_02561_),
    .B(_02564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08321_ (.Y(_02566_),
    .A(_02565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08322_ (.VDD(VPWR),
    .Y(_02567_),
    .A(\state[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08323_ (.Y(_02568_),
    .A(_02567_),
    .B(\state[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08324_ (.A(_02568_),
    .B(_02562_),
    .Y(_02569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout76 (.A(net93),
    .X(net76),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08326_ (.A(\state[2] ),
    .B(_02559_),
    .Y(_02571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08327_ (.A(\state[1] ),
    .B(_02567_),
    .Y(_02572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08328_ (.Y(_02573_),
    .A(_02571_),
    .B(_02572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08329_ (.VDD(VPWR),
    .Y(_02574_),
    .A(_02573_),
    .VSS(VGND));
 sg13g2_inv_1 _08330_ (.VDD(VPWR),
    .Y(_02575_),
    .A(_02568_),
    .VSS(VGND));
 sg13g2_nand2_2 _08331_ (.Y(_02576_),
    .A(_02575_),
    .B(_02571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1736 (.A(_04386_),
    .X(net1736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _08333_ (.A(_02576_),
    .Y(_02578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08334_ (.A(_02574_),
    .B(_02578_),
    .Y(_02579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08335_ (.VDD(VPWR),
    .Y(_02580_),
    .A(_02579_),
    .VSS(VGND));
 sg13g2_nor4_1 _08336_ (.A(_02563_),
    .B(_02566_),
    .C(_02569_),
    .D(_02580_),
    .Y(_02581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08337_ (.Y(_02582_),
    .A(\sipo.word_ready ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08338_ (.B(\sipo.word[10] ),
    .C(\sipo.word[9] ),
    .A(\sipo.word[11] ),
    .Y(_02583_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\sipo.word[8] ));
 sg13g2_nand4_1 _08339_ (.B(\sipo.word[14] ),
    .C(\sipo.word[13] ),
    .A(\sipo.word[15] ),
    .Y(_02584_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\sipo.word[12] ));
 sg13g2_nand4_1 _08340_ (.B(\sipo.word[2] ),
    .C(\sipo.word[1] ),
    .A(\sipo.word[3] ),
    .Y(_02585_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\sipo.word[0] ));
 sg13g2_nand4_1 _08341_ (.B(\sipo.word[6] ),
    .C(\sipo.word[5] ),
    .A(\sipo.word[7] ),
    .Y(_02586_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\sipo.word[4] ));
 sg13g2_nor4_1 _08342_ (.A(_02583_),
    .B(_02584_),
    .C(_02585_),
    .D(_02586_),
    .Y(_02587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08343_ (.A(_02582_),
    .B(_02576_),
    .C(_02587_),
    .Y(_00000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08344_ (.A(_02582_),
    .B(_02573_),
    .C(_02587_),
    .Y(_00001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08345_ (.A(_00000_),
    .B(_00001_),
    .Y(_02588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08346_ (.B1(_02588_),
    .VDD(VPWR),
    .Y(_02589_),
    .VSS(VGND),
    .A1(\sipo.word_ready ),
    .A2(_02581_));
 sg13g2_buf_1 place1716 (.A(_06574_),
    .X(net1716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08348_ (.Y(_02591_),
    .A(_02572_),
    .B(_02561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08349_ (.Y(_02592_),
    .A(_02591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08350_ (.Y(_02593_),
    .A(\instr[1] ),
    .B(\instr[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08351_ (.VDD(VPWR),
    .Y(_02594_),
    .A(_02593_),
    .VSS(VGND));
 sg13g2_nand2_1 _08352_ (.Y(_02595_),
    .A(_02592_),
    .B(_02594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _08353_ (.A(\instr[11] ),
    .B(\instr[10] ),
    .C(\instr[9] ),
    .D(\instr[8] ),
    .Y(_02596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _08354_ (.A(\instr[15] ),
    .B(\instr[14] ),
    .C(\instr[13] ),
    .D(\instr[12] ),
    .Y(_02597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08355_ (.Y(_02598_),
    .A(_02596_),
    .B(_02597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08356_ (.Y(_02599_),
    .A(_02598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _08357_ (.A(\instr[7] ),
    .B(\instr[6] ),
    .C(\instr[5] ),
    .Y(_02600_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\instr[4] ));
 sg13g2_inv_1 _08358_ (.VDD(VPWR),
    .Y(_02601_),
    .A(\instr[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08359_ (.A(\instr[3] ),
    .B(_02601_),
    .Y(_02602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08360_ (.B(_02600_),
    .C(_02602_),
    .A(_02599_),
    .Y(_02603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1737 (.A(net1736),
    .X(net1737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08362_ (.A(_02595_),
    .B(_02603_),
    .Y(_02605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08363_ (.VDD(VPWR),
    .Y(_02606_),
    .A(\instr[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08364_ (.A(\instr[1] ),
    .B(\instr[0] ),
    .Y(_02607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08365_ (.VDD(VPWR),
    .Y(_02608_),
    .A(_02607_),
    .VSS(VGND));
 sg13g2_nor3_1 _08366_ (.A(_02606_),
    .B(\instr[2] ),
    .C(_02608_),
    .Y(_02609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08367_ (.B(_02600_),
    .C(_02609_),
    .A(_02599_),
    .Y(_02610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08368_ (.A(\instr[3] ),
    .B(\instr[2] ),
    .Y(_02611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08369_ (.VDD(VPWR),
    .Y(_02612_),
    .A(\instr[0] ),
    .VSS(VGND));
 sg13g2_and3_1 _08370_ (.X(_02613_),
    .A(_02611_),
    .B(\instr[1] ),
    .C(_02612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08371_ (.B(_02600_),
    .C(_02613_),
    .A(_02599_),
    .Y(_02614_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08372_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02610_),
    .A2(_02614_),
    .Y(_02615_),
    .B1(_02591_));
 sg13g2_nor3_1 _08373_ (.A(_02605_),
    .B(_02615_),
    .C(_02589_),
    .Y(_02616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08374_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02559_),
    .A2(_02589_),
    .Y(_01361_),
    .B1(_02616_));
 sg13g2_nand4_1 _08375_ (.B(_02594_),
    .C(_02600_),
    .A(_02599_),
    .Y(_02617_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02611_));
 sg13g2_o21ai_1 _08376_ (.B1(_02617_),
    .VDD(VPWR),
    .Y(_02618_),
    .VSS(VGND),
    .A1(_02594_),
    .A2(_02603_));
 sg13g2_nand2_2 _08377_ (.Y(_02619_),
    .A(_02559_),
    .B(\state[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08378_ (.A(_02619_),
    .B_N(_02572_),
    .Y(_07115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08379_ (.Y(_02620_),
    .B(_07115_),
    .A_N(\fpdiv.reg2en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08380_ (.A(_02619_),
    .B_N(_02564_),
    .Y(_07116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08381_ (.Y(_02621_),
    .B(_07116_),
    .A_N(\fpmul.reg3en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08382_ (.A(_02568_),
    .B(_02619_),
    .Y(_07114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08383_ (.Y(_02622_),
    .B(_07114_),
    .A_N(\fp16_sum_pipe.reg4en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08384_ (.A(_02560_),
    .B(_02619_),
    .Y(_07113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08385_ (.VDD(VPWR),
    .Y(_02623_),
    .A(\fp16_res_pipe.reg4en.q[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08386_ (.Y(_02624_),
    .A(_07113_),
    .B(_02623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08387_ (.B(_02621_),
    .C(_02622_),
    .A(_02620_),
    .Y(_02625_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02624_));
 sg13g2_a21oi_1 _08388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02618_),
    .A2(_02563_),
    .Y(_02626_),
    .B1(_02625_));
 sg13g2_nor2_1 _08389_ (.A(_02626_),
    .B(_02589_),
    .Y(_01360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08390_ (.A(\instr[1] ),
    .B(_02612_),
    .Y(_02627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08391_ (.B(_02600_),
    .C(_02611_),
    .A(_02599_),
    .Y(_02628_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02627_));
 sg13g2_nand3b_1 _08392_ (.B(_02610_),
    .C(_02628_),
    .Y(_02629_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_02618_));
 sg13g2_o21ai_1 _08393_ (.B1(_02617_),
    .VDD(VPWR),
    .Y(_02630_),
    .VSS(VGND),
    .A1(_02608_),
    .A2(_02603_));
 sg13g2_nand2_1 _08394_ (.Y(_02631_),
    .A(_02630_),
    .B(_02563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout75 (.A(net76),
    .X(net75),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08396_ (.Y(_02633_),
    .A(_02618_),
    .B(_02569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08397_ (.B(_02633_),
    .C(_02622_),
    .A(_02631_),
    .Y(_02634_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02624_));
 sg13g2_a21oi_1 _08398_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02592_),
    .A2(_02629_),
    .Y(_02635_),
    .B1(_02634_));
 sg13g2_nand2_1 _08399_ (.Y(_02636_),
    .A(_02589_),
    .B(\state[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08400_ (.B1(_02636_),
    .VDD(VPWR),
    .Y(_01359_),
    .VSS(VGND),
    .A1(_02589_),
    .A2(_02635_));
 sg13g2_nand2_1 _08401_ (.Y(_02637_),
    .A(_02620_),
    .B(_02624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08402_ (.Y(_02638_),
    .A(_02563_),
    .B(_02612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08403_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02595_),
    .A2(_02638_),
    .Y(_02639_),
    .B1(_02603_));
 sg13g2_nor3_1 _08404_ (.A(_02566_),
    .B(_02637_),
    .C(_02639_),
    .Y(_02640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _08405_ (.A(_02640_),
    .B(_02633_),
    .X(_02641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08406_ (.Y(_02642_),
    .A(_02589_),
    .B(\state[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08407_ (.B1(_02642_),
    .VDD(VPWR),
    .Y(_01358_),
    .VSS(VGND),
    .A1(_02589_),
    .A2(_02641_));
 sg13g2_inv_1 _08408_ (.VDD(VPWR),
    .Y(_02643_),
    .A(\fpdiv.divider0.state ),
    .VSS(VGND));
 sg13g2_inv_2 _08409_ (.Y(_02644_),
    .A(\fpdiv.divider0.counter[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08410_ (.VDD(VPWR),
    .Y(_02645_),
    .A(\fpdiv.divider0.counter[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08411_ (.A(\fpdiv.divider0.counter[1] ),
    .B(\fpdiv.divider0.counter[0] ),
    .Y(_02646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08412_ (.VDD(VPWR),
    .Y(_02647_),
    .A(_02646_),
    .VSS(VGND));
 sg13g2_nor3_2 _08413_ (.A(_02644_),
    .B(_02645_),
    .C(_02647_),
    .Y(_02648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout78 (.A(net80),
    .X(net78),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08415_ (.A(_02643_),
    .B(_02648_),
    .Y(_02650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1731 (.A(net1730),
    .X(net1731),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08417_ (.A(_01756_),
    .B(_02650_),
    .Y(_02652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout124 (.A(net127),
    .X(net124),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _08419_ (.A(net1707),
    .Y(\fpdiv.divider0.en_r ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08420_ (.Y(_02654_),
    .A(_02650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1725 (.A(net1724),
    .X(net1725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08422_ (.VDD(VPWR),
    .Y(_02656_),
    .A(\fpdiv.divider0.remainder_reg[9] ),
    .VSS(VGND));
 sg13g2_inv_1 _08423_ (.VDD(VPWR),
    .Y(_02657_),
    .A(\fpdiv.divider0.remainder_reg[8] ),
    .VSS(VGND));
 sg13g2_inv_1 _08424_ (.VDD(VPWR),
    .Y(_02658_),
    .A(\fpdiv.divider0.remainder_reg[7] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _08425_ (.Y(_02659_),
    .A(\fpdiv.divider0.divisor_reg[6] ),
    .B(\fpdiv.divider0.remainder_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08426_ (.VDD(VPWR),
    .Y(_02660_),
    .A(_02659_),
    .VSS(VGND));
 sg13g2_xnor2_1 _08427_ (.Y(_02661_),
    .A(\fpdiv.divider0.divisor_reg[5] ),
    .B(\fpdiv.divider0.remainder_reg[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08428_ (.A(\fpdiv.divider0.remainder_reg[4] ),
    .B(_01774_),
    .Y(_02662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08429_ (.VDD(VPWR),
    .Y(_02663_),
    .A(_02662_),
    .VSS(VGND));
 sg13g2_nand2_1 _08430_ (.Y(_02664_),
    .A(_02661_),
    .B(_02663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08431_ (.VDD(VPWR),
    .Y(_02665_),
    .A(_02664_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08432_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01772_),
    .A2(\fpdiv.divider0.remainder_reg[5] ),
    .Y(_02666_),
    .B1(_02665_));
 sg13g2_nor2_1 _08433_ (.A(_02660_),
    .B(_02666_),
    .Y(_02667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _08434_ (.A2(\fpdiv.divider0.remainder_reg[6] ),
    .A1(_01770_),
    .B1(_02667_),
    .X(_02668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08435_ (.Y(_02669_),
    .A(\fpdiv.divider0.divisor_reg[7] ),
    .B(\fpdiv.divider0.remainder_reg[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08436_ (.Y(_02670_),
    .A(_02668_),
    .B(_02669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08437_ (.B1(_02670_),
    .VDD(VPWR),
    .Y(_02671_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.divisor_reg[7] ),
    .A2(_02658_));
 sg13g2_xnor2_1 _08438_ (.Y(_02672_),
    .A(\fpdiv.divider0.divisor_reg[8] ),
    .B(\fpdiv.divider0.remainder_reg[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08439_ (.Y(_02673_),
    .A(_02671_),
    .B(_02672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08440_ (.B1(_02673_),
    .VDD(VPWR),
    .Y(_02674_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.divisor_reg[8] ),
    .A2(_02657_));
 sg13g2_xnor2_1 _08441_ (.Y(_02675_),
    .A(\fpdiv.divider0.divisor_reg[9] ),
    .B(\fpdiv.divider0.remainder_reg[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08442_ (.Y(_02676_),
    .A(_02674_),
    .B(_02675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08443_ (.B1(_02676_),
    .VDD(VPWR),
    .Y(_02677_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.divisor_reg[9] ),
    .A2(_02656_));
 sg13g2_xnor2_1 _08444_ (.Y(_02678_),
    .A(\fpdiv.divider0.divisor_reg[10] ),
    .B(\fpdiv.divider0.remainder_reg[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08445_ (.Y(_02679_),
    .A(_02677_),
    .B(_02678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08446_ (.Y(_02680_),
    .A(_01760_),
    .B(\fpdiv.divider0.remainder_reg[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08447_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02679_),
    .A2(_02680_),
    .Y(_02681_),
    .B1(\fpdiv.divider0.divisor_reg[11] ));
 sg13g2_and3_1 _08448_ (.X(_02682_),
    .A(_02679_),
    .B(\fpdiv.divider0.divisor_reg[11] ),
    .C(_02680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08449_ (.A(_02681_),
    .B(_02682_),
    .Y(_02683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08450_ (.VDD(VPWR),
    .Y(_02684_),
    .A(\fpdiv.divider0.remainder_reg[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08451_ (.Y(_02685_),
    .A(_02683_),
    .B(_02684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08452_ (.B1(_02685_),
    .VDD(VPWR),
    .Y(_02686_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.remainder_reg[11] ),
    .A2(_02683_));
 sg13g2_buf_2 fanout123 (.A(net124),
    .X(net123),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08454_ (.Y(_02688_),
    .A(_02652_),
    .B(\fpdiv.divider0.remainder_reg[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08455_ (.B1(_02688_),
    .VDD(VPWR),
    .Y(_01357_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02686_));
 sg13g2_inv_1 _08456_ (.VDD(VPWR),
    .Y(_02689_),
    .A(\fpdiv.divider0.remainder_reg[11] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08457_ (.A(\fpdiv.divider0.remainder_reg[11] ),
    .B(_02681_),
    .Y(_02690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08458_ (.A(_02682_),
    .B(_02690_),
    .Y(_02691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08459_ (.Y(_02692_),
    .A(_02684_),
    .B(_02691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_92_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_92_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_91_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_91_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _08462_ (.B(_02677_),
    .A(_02678_),
    .X(_02695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08463_ (.A(net1647),
    .B_N(\fpdiv.divider0.remainder_reg[10] ),
    .Y(_02696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08464_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1647),
    .A2(_02695_),
    .Y(_02697_),
    .B1(_02696_));
 sg13g2_a22oi_1 _08465_ (.Y(_01356_),
    .B1(net1718),
    .B2(_02697_),
    .A2(_02652_),
    .A1(_02689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08466_ (.Y(_02698_),
    .A(_02675_),
    .B(_02674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08467_ (.Y(_02699_),
    .A(net1647),
    .B(_02698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08468_ (.B1(_02699_),
    .VDD(VPWR),
    .Y(_02700_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.remainder_reg[9] ),
    .A2(net1647));
 sg13g2_a22oi_1 _08469_ (.Y(_02701_),
    .B1(\fpdiv.divider0.remainder_reg[10] ),
    .B2(net1708),
    .A2(_01756_),
    .A1(\fpdiv.divider0.dividend[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08470_ (.B1(_02701_),
    .VDD(VPWR),
    .Y(_01355_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02700_));
 sg13g2_xnor2_1 _08471_ (.Y(_02702_),
    .A(_02672_),
    .B(_02671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08472_ (.Y(_02703_),
    .A(net1647),
    .B(_02702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08473_ (.B1(_02703_),
    .VDD(VPWR),
    .Y(_02704_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.remainder_reg[8] ),
    .A2(net1647));
 sg13g2_a22oi_1 _08474_ (.Y(_02705_),
    .B1(\fpdiv.divider0.remainder_reg[9] ),
    .B2(net1708),
    .A2(_01756_),
    .A1(\fpdiv.divider0.dividend[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08475_ (.B1(_02705_),
    .VDD(VPWR),
    .Y(_01354_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02704_));
 sg13g2_xnor2_1 _08476_ (.Y(_02706_),
    .A(_02669_),
    .B(_02668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08477_ (.Y(_02707_),
    .A(_02692_),
    .B(_02706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08478_ (.B1(_02707_),
    .VDD(VPWR),
    .Y(_02708_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.remainder_reg[7] ),
    .A2(net1647));
 sg13g2_a22oi_1 _08479_ (.Y(_02709_),
    .B1(\fpdiv.divider0.remainder_reg[8] ),
    .B2(net1708),
    .A2(net1748),
    .A1(\fpdiv.divider0.dividend[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08480_ (.B1(_02709_),
    .VDD(VPWR),
    .Y(_01353_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02708_));
 sg13g2_nand2_1 _08481_ (.Y(_02710_),
    .A(_02666_),
    .B(_02660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08482_ (.VDD(VPWR),
    .Y(_02711_),
    .A(_02710_),
    .VSS(VGND));
 sg13g2_o21ai_1 _08483_ (.B1(_02692_),
    .VDD(VPWR),
    .Y(_02712_),
    .VSS(VGND),
    .A1(_02667_),
    .A2(_02711_));
 sg13g2_o21ai_1 _08484_ (.B1(_02712_),
    .VDD(VPWR),
    .Y(_02713_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.remainder_reg[6] ),
    .A2(_02692_));
 sg13g2_a22oi_1 _08485_ (.Y(_02714_),
    .B1(\fpdiv.divider0.remainder_reg[7] ),
    .B2(net1708),
    .A2(net1748),
    .A1(\fpdiv.divider0.dividend[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08486_ (.B1(_02714_),
    .VDD(VPWR),
    .Y(_01352_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02713_));
 sg13g2_nor2_1 _08487_ (.A(_02663_),
    .B(_02661_),
    .Y(_02715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08488_ (.B1(_02692_),
    .VDD(VPWR),
    .Y(_02716_),
    .VSS(VGND),
    .A1(_02665_),
    .A2(_02715_));
 sg13g2_o21ai_1 _08489_ (.B1(_02716_),
    .VDD(VPWR),
    .Y(_02717_),
    .VSS(VGND),
    .A1(\fpdiv.divider0.remainder_reg[5] ),
    .A2(_02692_));
 sg13g2_a22oi_1 _08490_ (.Y(_02718_),
    .B1(\fpdiv.divider0.remainder_reg[6] ),
    .B2(net1708),
    .A2(net1748),
    .A1(\fpdiv.divider0.dividend[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08491_ (.B1(_02718_),
    .VDD(VPWR),
    .Y(_01351_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02717_));
 sg13g2_nand2_1 _08492_ (.Y(_02719_),
    .A(_02692_),
    .B(\fpdiv.divider0.divisor_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _08493_ (.B(_02719_),
    .A(\fpdiv.divider0.remainder_reg[4] ),
    .X(_02720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08494_ (.Y(_02721_),
    .B1(\fpdiv.divider0.remainder_reg[5] ),
    .B2(net1708),
    .A2(net1748),
    .A1(\fpdiv.divider0.dividend[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08495_ (.B1(_02721_),
    .VDD(VPWR),
    .Y(_01350_),
    .VSS(VGND),
    .A1(net1705),
    .A2(_02720_));
 sg13g2_inv_2 _08496_ (.Y(_02722_),
    .A(\fpdiv.divider0.dividend[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08497_ (.Y(_02723_),
    .A(net1708),
    .B(\fpdiv.divider0.remainder_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08498_ (.B1(_02723_),
    .VDD(VPWR),
    .Y(_01349_),
    .VSS(VGND),
    .A1(_02722_),
    .A2(_01758_));
 sg13g2_xor2_1 _08499_ (.B(\acc_sum.op_sign_logic0.s_b ),
    .A(\acc_sum.op_sign_logic0.s_a ),
    .X(_02724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1851 (.A(\fpdiv.div_out[11] ),
    .X(net1851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08501_ (.VDD(VPWR),
    .Y(_02726_),
    .A(_02724_),
    .VSS(VGND));
 sg13g2_buf_2 fanout79 (.A(net80),
    .X(net79),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08503_ (.A(\acc_sum.seg_reg1.q[21] ),
    .B(net1816),
    .Y(_02728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08504_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1740),
    .A2(net1816),
    .Y(_01348_),
    .B1(_02728_));
 sg13g2_inv_1 _08505_ (.VDD(VPWR),
    .Y(_02729_),
    .A(\acc_sum.seg_reg1.q[20] ),
    .VSS(VGND));
 sg13g2_nor2b_1 _08506_ (.A(\acc_sum.op_sign_logic0.mantisa_a[9] ),
    .B_N(\acc_sum.op_sign_logic0.mantisa_b[9] ),
    .Y(_02730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08507_ (.A(\acc_sum.op_sign_logic0.mantisa_b[9] ),
    .B_N(\acc_sum.op_sign_logic0.mantisa_a[9] ),
    .Y(_02731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08508_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08509_ (.A(\acc_sum.op_sign_logic0.mantisa_a[8] ),
    .B_N(\acc_sum.op_sign_logic0.mantisa_b[8] ),
    .Y(_02733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08510_ (.VDD(VPWR),
    .Y(_02734_),
    .A(\acc_sum.op_sign_logic0.mantisa_b[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08511_ (.A(\acc_sum.op_sign_logic0.mantisa_a[7] ),
    .B(_02734_),
    .Y(_02735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08512_ (.A(\acc_sum.op_sign_logic0.mantisa_b[7] ),
    .B_N(\acc_sum.op_sign_logic0.mantisa_a[7] ),
    .Y(_02736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08513_ (.A(_02735_),
    .B(_02736_),
    .Y(_02737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08514_ (.VDD(VPWR),
    .Y(_02738_),
    .A(_02737_),
    .VSS(VGND));
 sg13g2_inv_1 _08515_ (.VDD(VPWR),
    .Y(_02739_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[6] ),
    .VSS(VGND));
 sg13g2_nor2_2 _08516_ (.A(\acc_sum.op_sign_logic0.mantisa_b[6] ),
    .B(_02739_),
    .Y(_02740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08517_ (.Y(_02741_),
    .A(_02739_),
    .B(\acc_sum.op_sign_logic0.mantisa_b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08518_ (.VDD(VPWR),
    .Y(_02742_),
    .A(_02741_),
    .VSS(VGND));
 sg13g2_nor2_1 _08519_ (.A(_02740_),
    .B(_02742_),
    .Y(_02743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08520_ (.VDD(VPWR),
    .Y(_02744_),
    .A(_02743_),
    .VSS(VGND));
 sg13g2_nor2_1 _08521_ (.A(_02738_),
    .B(_02744_),
    .Y(_02745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08522_ (.VDD(VPWR),
    .Y(_02746_),
    .A(_02745_),
    .VSS(VGND));
 sg13g2_inv_1 _08523_ (.VDD(VPWR),
    .Y(_02747_),
    .A(\acc_sum.op_sign_logic0.mantisa_b[2] ),
    .VSS(VGND));
 sg13g2_nor2_2 _08524_ (.A(\acc_sum.op_sign_logic0.mantisa_a[2] ),
    .B(_02747_),
    .Y(_02748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08525_ (.VDD(VPWR),
    .Y(_02749_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08526_ (.A(\acc_sum.op_sign_logic0.mantisa_b[3] ),
    .B(_02749_),
    .Y(_02750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08527_ (.Y(_02751_),
    .A(_02749_),
    .B(\acc_sum.op_sign_logic0.mantisa_b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08528_ (.VDD(VPWR),
    .Y(_02752_),
    .A(_02751_),
    .VSS(VGND));
 sg13g2_nor2_1 _08529_ (.A(_02750_),
    .B(_02752_),
    .Y(_02753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08530_ (.Y(_02754_),
    .A(_02747_),
    .B(\acc_sum.op_sign_logic0.mantisa_a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08531_ (.VDD(VPWR),
    .Y(_02755_),
    .A(_02754_),
    .VSS(VGND));
 sg13g2_nor2_2 _08532_ (.A(_02748_),
    .B(_02755_),
    .Y(_02756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08533_ (.VDD(VPWR),
    .Y(_02757_),
    .A(_02756_),
    .VSS(VGND));
 sg13g2_inv_1 _08534_ (.VDD(VPWR),
    .Y(_02758_),
    .A(_02753_),
    .VSS(VGND));
 sg13g2_nor2_1 _08535_ (.A(_02757_),
    .B(_02758_),
    .Y(_02759_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _08536_ (.Y(_02760_),
    .B(\acc_sum.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\acc_sum.op_sign_logic0.mantisa_b[1] ));
 sg13g2_inv_1 _08537_ (.VDD(VPWR),
    .Y(_02761_),
    .A(\acc_sum.op_sign_logic0.mantisa_b[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08538_ (.Y(_02762_),
    .A(_02761_),
    .B(\acc_sum.op_sign_logic0.mantisa_a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08539_ (.VDD(VPWR),
    .Y(_02763_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08540_ (.Y(_02764_),
    .A(_02763_),
    .B(\acc_sum.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08541_ (.VDD(VPWR),
    .Y(_02765_),
    .A(_02764_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08542_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02760_),
    .A2(_02762_),
    .Y(_02766_),
    .B1(_02765_));
 sg13g2_inv_1 _08543_ (.VDD(VPWR),
    .Y(_02767_),
    .A(_02766_),
    .VSS(VGND));
 sg13g2_a221oi_1 _08544_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02767_),
    .C1(_02752_),
    .B1(_02759_),
    .A1(_02748_),
    .Y(_02768_),
    .A2(_02753_));
 sg13g2_inv_1 _08545_ (.VDD(VPWR),
    .Y(_02769_),
    .A(_02768_),
    .VSS(VGND));
 sg13g2_inv_1 _08546_ (.VDD(VPWR),
    .Y(_02770_),
    .A(\acc_sum.op_sign_logic0.mantisa_b[4] ),
    .VSS(VGND));
 sg13g2_nor2_2 _08547_ (.A(\acc_sum.op_sign_logic0.mantisa_a[4] ),
    .B(_02770_),
    .Y(_02771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08548_ (.Y(_02772_),
    .A(_02770_),
    .B(\acc_sum.op_sign_logic0.mantisa_a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08549_ (.VDD(VPWR),
    .Y(_02773_),
    .A(_02772_),
    .VSS(VGND));
 sg13g2_nor2_2 _08550_ (.A(_02771_),
    .B(_02773_),
    .Y(_02774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08551_ (.VDD(VPWR),
    .Y(_02775_),
    .A(_02774_),
    .VSS(VGND));
 sg13g2_inv_1 _08552_ (.VDD(VPWR),
    .Y(_02776_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08553_ (.A(\acc_sum.op_sign_logic0.mantisa_b[5] ),
    .B(_02776_),
    .Y(_02777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08554_ (.Y(_02778_),
    .A(_02776_),
    .B(\acc_sum.op_sign_logic0.mantisa_b[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08555_ (.VDD(VPWR),
    .Y(_02779_),
    .A(_02778_),
    .VSS(VGND));
 sg13g2_nor2_1 _08556_ (.A(_02777_),
    .B(_02779_),
    .Y(_02780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08557_ (.VDD(VPWR),
    .Y(_02781_),
    .A(_02780_),
    .VSS(VGND));
 sg13g2_nor2_1 _08558_ (.A(_02775_),
    .B(_02781_),
    .Y(_02782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08559_ (.VDD(VPWR),
    .Y(_02783_),
    .A(_02771_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08560_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02783_),
    .A2(_02778_),
    .Y(_02784_),
    .B1(_02777_));
 sg13g2_a21oi_1 _08561_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02769_),
    .A2(_02782_),
    .Y(_02785_),
    .B1(_02784_));
 sg13g2_a21oi_1 _08562_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02737_),
    .A2(_02742_),
    .Y(_02786_),
    .B1(_02735_));
 sg13g2_o21ai_1 _08563_ (.B1(_02786_),
    .VDD(VPWR),
    .Y(_02787_),
    .VSS(VGND),
    .A1(_02746_),
    .A2(_02785_));
 sg13g2_inv_2 _08564_ (.Y(_02788_),
    .A(_02732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08565_ (.A(\acc_sum.op_sign_logic0.mantisa_b[8] ),
    .B_N(\acc_sum.op_sign_logic0.mantisa_a[8] ),
    .Y(_02789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08566_ (.A(_02789_),
    .B(_02733_),
    .Y(_02790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08567_ (.VDD(VPWR),
    .Y(_02791_),
    .A(_02790_),
    .VSS(VGND));
 sg13g2_nor2_1 _08568_ (.A(_02788_),
    .B(_02791_),
    .Y(_02792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _08569_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02792_),
    .C1(_02730_),
    .B1(_02787_),
    .A1(_02732_),
    .Y(_02793_),
    .A2(_02733_));
 sg13g2_inv_1 _08570_ (.VDD(VPWR),
    .Y(_02794_),
    .A(_02793_),
    .VSS(VGND));
 sg13g2_inv_1 _08571_ (.VDD(VPWR),
    .Y(_02795_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08572_ (.A(\acc_sum.op_sign_logic0.mantisa_b[10] ),
    .B(_02795_),
    .Y(_02796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08573_ (.VDD(VPWR),
    .Y(_02797_),
    .A(\acc_sum.op_sign_logic0.mantisa_b[10] ),
    .VSS(VGND));
 sg13g2_nor2_2 _08574_ (.A(\acc_sum.op_sign_logic0.mantisa_a[10] ),
    .B(_02797_),
    .Y(_02798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08575_ (.A(_02796_),
    .B(_02798_),
    .Y(_02799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08576_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_02798_),
    .Y(_02800_),
    .A2(_02799_),
    .A1(_02794_));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08578_ (.VDD(VPWR),
    .Y(_02802_),
    .A(\acc_sum.op_sign_logic0.s_a ),
    .VSS(VGND));
 sg13g2_inv_2 _08579_ (.Y(_02803_),
    .A(\acc_sum.reg2en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08580_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02800_),
    .A2(_02802_),
    .Y(_02804_),
    .B1(_02803_));
 sg13g2_o21ai_1 _08581_ (.B1(_02804_),
    .VDD(VPWR),
    .Y(_02805_),
    .VSS(VGND),
    .A1(\acc_sum.op_sign_logic0.s_b ),
    .A2(_02800_));
 sg13g2_o21ai_1 _08582_ (.B1(_02805_),
    .VDD(VPWR),
    .Y(_01347_),
    .VSS(VGND),
    .A1(net1814),
    .A2(_02729_));
 sg13g2_inv_4 _08583_ (.A(\acc_sum.add_renorm0.mantisa[11] ),
    .Y(_02806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08584_ (.Y(_02807_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[10] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08585_ (.B1(\acc_sum.reg2en.q[0] ),
    .VDD(VPWR),
    .Y(_02808_),
    .VSS(VGND),
    .A1(_02807_),
    .A2(_02724_));
 sg13g2_nand2_1 _08586_ (.Y(_02809_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[9] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08587_ (.VDD(VPWR),
    .Y(_02810_),
    .A(_02809_),
    .VSS(VGND));
 sg13g2_nand2_1 _08588_ (.Y(_02811_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[8] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08589_ (.A(_02811_),
    .B(_02724_),
    .Y(_02812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08590_ (.A(\acc_sum.op_sign_logic0.mantisa_a[7] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[7] ),
    .Y(_02813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08591_ (.Y(_02814_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[6] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08592_ (.VDD(VPWR),
    .Y(_02815_),
    .A(_02814_),
    .VSS(VGND));
 sg13g2_nand2_2 _08593_ (.Y(_02816_),
    .A(_02760_),
    .B(_02764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08594_ (.Y(_02817_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[0] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08595_ (.VDD(VPWR),
    .Y(_02818_),
    .A(_02817_),
    .VSS(VGND));
 sg13g2_nand2_1 _08596_ (.Y(_02819_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[1] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08597_ (.VDD(VPWR),
    .Y(_02820_),
    .A(_02819_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08598_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02816_),
    .A2(_02818_),
    .Y(_02821_),
    .B1(_02820_));
 sg13g2_nand2_1 _08599_ (.Y(_02822_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[2] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08600_ (.B1(_02822_),
    .VDD(VPWR),
    .Y(_02823_),
    .VSS(VGND),
    .A1(_02756_),
    .A2(_02821_));
 sg13g2_nand2_1 _08601_ (.Y(_02824_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[3] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08602_ (.VDD(VPWR),
    .Y(_02825_),
    .A(_02824_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02823_),
    .A2(_02758_),
    .Y(_02826_),
    .B1(_02825_));
 sg13g2_nand2_1 _08604_ (.Y(_02827_),
    .A(\acc_sum.op_sign_logic0.mantisa_a[4] ),
    .B(\acc_sum.op_sign_logic0.mantisa_b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08605_ (.B1(_02827_),
    .VDD(VPWR),
    .Y(_02828_),
    .VSS(VGND),
    .A1(_02774_),
    .A2(_02826_));
 sg13g2_nand2_1 _08606_ (.Y(_02829_),
    .A(_02828_),
    .B(net1739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08607_ (.B(\acc_sum.op_sign_logic0.mantisa_a[5] ),
    .C(\acc_sum.op_sign_logic0.mantisa_b[5] ),
    .A(net1739),
    .Y(_02830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08608_ (.B1(_02830_),
    .VDD(VPWR),
    .Y(_02831_),
    .VSS(VGND),
    .A1(_02780_),
    .A2(_02829_));
 sg13g2_a22oi_1 _08609_ (.Y(_02832_),
    .B1(_02744_),
    .B2(_02831_),
    .A2(_02815_),
    .A1(_02726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08610_ (.B(\acc_sum.op_sign_logic0.mantisa_a[7] ),
    .C(\acc_sum.op_sign_logic0.mantisa_b[7] ),
    .A(net1740),
    .Y(_02833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08611_ (.B1(_02833_),
    .VDD(VPWR),
    .Y(_02834_),
    .VSS(VGND),
    .A1(_02813_),
    .A2(_02832_));
 sg13g2_nand2_1 _08612_ (.Y(_02835_),
    .A(_02834_),
    .B(_02791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08613_ (.Y(_02836_),
    .B(_02835_),
    .A_N(_02812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08614_ (.Y(_02837_),
    .B1(_02788_),
    .B2(_02836_),
    .A2(_02810_),
    .A1(net1740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08615_ (.A(_02799_),
    .B(_02837_),
    .Y(_02838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08616_ (.A(_02808_),
    .B(_02838_),
    .Y(_02839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02803_),
    .A2(_02806_),
    .Y(_01346_),
    .B1(_02839_));
 sg13g2_inv_1 _08618_ (.VDD(VPWR),
    .Y(_02840_),
    .A(_02799_),
    .VSS(VGND));
 sg13g2_nor2_2 _08619_ (.A(\acc_sum.op_sign_logic0.mantisa_a[0] ),
    .B(_02761_),
    .Y(_02841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08620_ (.VDD(VPWR),
    .Y(_02842_),
    .A(_02762_),
    .VSS(VGND));
 sg13g2_nor4_1 _08621_ (.A(_02841_),
    .B(_02842_),
    .C(_02816_),
    .D(_02840_),
    .Y(_02843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _08622_ (.A(_02792_),
    .B(_02759_),
    .C(_02782_),
    .D(_02745_),
    .X(_02844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08623_ (.B1(_02760_),
    .VDD(VPWR),
    .Y(_02845_),
    .VSS(VGND),
    .A1(_02841_),
    .A2(_02765_));
 sg13g2_a21oi_1 _08624_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02845_),
    .A2(_02756_),
    .Y(_02846_),
    .B1(_02755_));
 sg13g2_inv_1 _08625_ (.VDD(VPWR),
    .Y(_02847_),
    .A(_02846_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08626_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02847_),
    .A2(_02751_),
    .Y(_02848_),
    .B1(_02750_));
 sg13g2_inv_1 _08627_ (.VDD(VPWR),
    .Y(_02849_),
    .A(_02848_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02849_),
    .A2(_02774_),
    .Y(_02850_),
    .B1(_02773_));
 sg13g2_inv_1 _08629_ (.VDD(VPWR),
    .Y(_02851_),
    .A(_02850_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02851_),
    .A2(_02778_),
    .Y(_02852_),
    .B1(_02777_));
 sg13g2_a21oi_1 _08631_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02737_),
    .A2(_02740_),
    .Y(_02853_),
    .B1(_02736_));
 sg13g2_o21ai_1 _08632_ (.B1(_02853_),
    .VDD(VPWR),
    .Y(_02854_),
    .VSS(VGND),
    .A1(_02746_),
    .A2(_02852_));
 sg13g2_nand2_1 _08633_ (.Y(_02855_),
    .A(_02854_),
    .B(_02792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08634_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02732_),
    .A2(_02789_),
    .Y(_02856_),
    .B1(_02731_));
 sg13g2_a221oi_1 _08635_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02856_),
    .C1(_02798_),
    .B1(_02855_),
    .A1(_02843_),
    .Y(_02857_),
    .A2(_02844_));
 sg13g2_o21ai_1 _08636_ (.B1(_02724_),
    .VDD(VPWR),
    .Y(_02858_),
    .VSS(VGND),
    .A1(_02796_),
    .A2(_02793_));
 sg13g2_o21ai_1 _08637_ (.B1(_02837_),
    .VDD(VPWR),
    .Y(_02859_),
    .VSS(VGND),
    .A1(_02857_),
    .A2(_02858_));
 sg13g2_xnor2_1 _08638_ (.Y(_02860_),
    .A(_02840_),
    .B(_02859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08639_ (.A(net1818),
    .B(\acc_sum.add_renorm0.mantisa[10] ),
    .Y(_02861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08640_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02860_),
    .A2(net1818),
    .Y(_01345_),
    .B1(_02861_));
 sg13g2_a21oi_1 _08641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02787_),
    .A2(_02790_),
    .Y(_02862_),
    .B1(_02733_));
 sg13g2_nor2_1 _08642_ (.A(_02862_),
    .B(net1671),
    .Y(_02863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08643_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02854_),
    .A2(_02790_),
    .Y(_02864_),
    .B1(_02789_));
 sg13g2_inv_1 _08644_ (.VDD(VPWR),
    .Y(_02865_),
    .A(_02800_),
    .VSS(VGND));
 sg13g2_o21ai_1 _08645_ (.B1(_02724_),
    .VDD(VPWR),
    .Y(_02866_),
    .VSS(VGND),
    .A1(_02864_),
    .A2(_02865_));
 sg13g2_inv_1 _08646_ (.VDD(VPWR),
    .Y(_02867_),
    .A(_02836_),
    .VSS(VGND));
 sg13g2_o21ai_1 _08647_ (.B1(_02867_),
    .VDD(VPWR),
    .Y(_02868_),
    .VSS(VGND),
    .A1(_02863_),
    .A2(_02866_));
 sg13g2_xnor2_1 _08648_ (.Y(_02869_),
    .A(_02788_),
    .B(_02868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08649_ (.A(net1816),
    .B(\acc_sum.add_renorm0.mantisa[9] ),
    .Y(_02870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08650_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02869_),
    .A2(net1816),
    .Y(_01344_),
    .B1(_02870_));
 sg13g2_a21oi_1 _08651_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1671),
    .A2(_02854_),
    .Y(_02871_),
    .B1(net1740));
 sg13g2_nand2_1 _08652_ (.Y(_02872_),
    .A(_02865_),
    .B(_02787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02871_),
    .A2(_02872_),
    .Y(_02873_),
    .B1(_02834_));
 sg13g2_xnor2_1 _08654_ (.Y(_02874_),
    .A(_02790_),
    .B(_02873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08655_ (.A(net1818),
    .B(\acc_sum.add_renorm0.mantisa[8] ),
    .Y(_02875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08656_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02874_),
    .A2(net1818),
    .Y(_01343_),
    .B1(_02875_));
 sg13g2_inv_1 _08657_ (.VDD(VPWR),
    .Y(_02876_),
    .A(_02852_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02876_),
    .A2(_02743_),
    .Y(_02877_),
    .B1(_02740_));
 sg13g2_a21oi_1 _08659_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02785_),
    .A2(_02741_),
    .Y(_02878_),
    .B1(_02740_));
 sg13g2_nand2_1 _08660_ (.Y(_02879_),
    .A(net1668),
    .B(_02878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08661_ (.B1(_02879_),
    .VDD(VPWR),
    .Y(_02880_),
    .VSS(VGND),
    .A1(net1668),
    .A2(_02877_));
 sg13g2_o21ai_1 _08662_ (.B1(_02832_),
    .VDD(VPWR),
    .Y(_02881_),
    .VSS(VGND),
    .A1(net1740),
    .A2(_02880_));
 sg13g2_xnor2_1 _08663_ (.Y(_02882_),
    .A(_02738_),
    .B(_02881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08664_ (.A(net1818),
    .B(\acc_sum.add_renorm0.mantisa[7] ),
    .Y(_02883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08665_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02882_),
    .A2(net1818),
    .Y(_01342_),
    .B1(_02883_));
 sg13g2_a21oi_1 _08666_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1671),
    .A2(_02876_),
    .Y(_02884_),
    .B1(net1740));
 sg13g2_nand2b_1 _08667_ (.Y(_02885_),
    .B(net1668),
    .A_N(_02785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02884_),
    .A2(_02885_),
    .Y(_02886_),
    .B1(_02831_));
 sg13g2_xnor2_1 _08669_ (.Y(_02887_),
    .A(_02743_),
    .B(_02886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08670_ (.A(net1818),
    .B(\acc_sum.add_renorm0.mantisa[6] ),
    .Y(_02888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08671_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02887_),
    .A2(net1818),
    .Y(_01341_),
    .B1(_02888_));
 sg13g2_a21oi_1 _08672_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02769_),
    .A2(_02774_),
    .Y(_02889_),
    .B1(_02771_));
 sg13g2_nor2_1 _08673_ (.A(_02889_),
    .B(net1671),
    .Y(_02890_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08674_ (.B1(_02724_),
    .VDD(VPWR),
    .Y(_02891_),
    .VSS(VGND),
    .A1(_02850_),
    .A2(net1668));
 sg13g2_o21ai_1 _08675_ (.B1(_02829_),
    .VDD(VPWR),
    .Y(_02892_),
    .VSS(VGND),
    .A1(_02890_),
    .A2(_02891_));
 sg13g2_xnor2_1 _08676_ (.Y(_02893_),
    .A(_02781_),
    .B(_02892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08677_ (.A(net1816),
    .B(\acc_sum.add_renorm0.mantisa[5] ),
    .Y(_02894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08678_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02893_),
    .A2(net1816),
    .Y(_01340_),
    .B1(_02894_));
 sg13g2_inv_1 _08679_ (.VDD(VPWR),
    .Y(_02895_),
    .A(_02826_),
    .VSS(VGND));
 sg13g2_nand2_1 _08680_ (.Y(_02896_),
    .A(net1668),
    .B(_02769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08681_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1671),
    .A2(_02849_),
    .Y(_02897_),
    .B1(net1739));
 sg13g2_a22oi_1 _08682_ (.Y(_02898_),
    .B1(_02896_),
    .B2(_02897_),
    .A2(_02895_),
    .A1(net1739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08683_ (.Y(_02899_),
    .A(_02774_),
    .B(_02898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08684_ (.A(net1817),
    .B(\acc_sum.add_renorm0.mantisa[4] ),
    .Y(_02900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08685_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02899_),
    .A2(net1817),
    .Y(_01339_),
    .B1(_02900_));
 sg13g2_nor2_1 _08686_ (.A(_02757_),
    .B(_02766_),
    .Y(_02901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08687_ (.B1(net1668),
    .VDD(VPWR),
    .Y(_02902_),
    .VSS(VGND),
    .A1(_02748_),
    .A2(_02901_));
 sg13g2_a21oi_1 _08688_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1671),
    .A2(_02847_),
    .Y(_02903_),
    .B1(net1739));
 sg13g2_a22oi_1 _08689_ (.Y(_02904_),
    .B1(_02902_),
    .B2(_02903_),
    .A2(_02823_),
    .A1(net1739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08690_ (.Y(_02905_),
    .A(_02753_),
    .B(_02904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08691_ (.A(net1817),
    .B(\acc_sum.add_renorm0.mantisa[3] ),
    .Y(_02906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08692_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02905_),
    .A2(net1817),
    .Y(_01338_),
    .B1(_02906_));
 sg13g2_inv_1 _08693_ (.VDD(VPWR),
    .Y(_02907_),
    .A(_02821_),
    .VSS(VGND));
 sg13g2_nand2_1 _08694_ (.Y(_02908_),
    .A(net1668),
    .B(_02767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08695_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1671),
    .A2(_02845_),
    .Y(_02909_),
    .B1(net1739));
 sg13g2_a22oi_1 _08696_ (.Y(_02910_),
    .B1(_02908_),
    .B2(_02909_),
    .A2(_02907_),
    .A1(net1739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08697_ (.Y(_02911_),
    .A(_02756_),
    .B(_02910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08698_ (.A(net1817),
    .B(\acc_sum.add_renorm0.mantisa[2] ),
    .Y(_02912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08699_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02911_),
    .A2(net1817),
    .Y(_01337_),
    .B1(_02912_));
 sg13g2_nand2_1 _08700_ (.Y(_02913_),
    .A(net1668),
    .B(_02842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1671),
    .A2(_02841_),
    .Y(_02914_),
    .B1(net1740));
 sg13g2_a22oi_1 _08702_ (.Y(_02915_),
    .B1(_02913_),
    .B2(_02914_),
    .A2(_02817_),
    .A1(net1740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08703_ (.Y(_02916_),
    .A(_02816_),
    .B(_02915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08704_ (.A(net1817),
    .B(\acc_sum.add_renorm0.mantisa[1] ),
    .Y(_02917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08705_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02916_),
    .A2(net1817),
    .Y(_01336_),
    .B1(_02917_));
 sg13g2_inv_1 _08706_ (.VDD(VPWR),
    .Y(_02918_),
    .A(\acc_sum.add_renorm0.mantisa[0] ),
    .VSS(VGND));
 sg13g2_nor3_1 _08707_ (.A(_02803_),
    .B(_02841_),
    .C(_02842_),
    .Y(_02919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08708_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02803_),
    .A2(_02918_),
    .Y(_01335_),
    .B1(_02919_));
 sg13g2_inv_2 _08709_ (.Y(_02920_),
    .A(\acc_sum.add_renorm0.exp[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08710_ (.Y(_02921_),
    .A(net1819),
    .B(\acc_sum.seg_reg0.q[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08711_ (.B1(_02921_),
    .VDD(VPWR),
    .Y(_01334_),
    .VSS(VGND),
    .A1(net1814),
    .A2(_02920_));
 sg13g2_inv_1 _08712_ (.VDD(VPWR),
    .Y(_02922_),
    .A(\acc_sum.seg_reg0.q[28] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08713_ (.A(net1814),
    .B(\acc_sum.add_renorm0.exp[6] ),
    .Y(_02923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08714_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1814),
    .A2(_02922_),
    .Y(_01333_),
    .B1(_02923_));
 sg13g2_inv_2 _08715_ (.Y(_02924_),
    .A(\acc_sum.add_renorm0.exp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08716_ (.Y(_02925_),
    .A(net1819),
    .B(\acc_sum.seg_reg0.q[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08717_ (.B1(_02925_),
    .VDD(VPWR),
    .Y(_01332_),
    .VSS(VGND),
    .A1(net1814),
    .A2(_02924_));
 sg13g2_mux2_1 _08718_ (.A0(\acc_sum.add_renorm0.exp[4] ),
    .A1(\acc_sum.seg_reg0.q[26] ),
    .S(net1819),
    .X(_01331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08719_ (.VDD(VPWR),
    .Y(_02926_),
    .A(\acc_sum.add_renorm0.exp[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08720_ (.Y(_02927_),
    .A(net1819),
    .B(\acc_sum.seg_reg0.q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08721_ (.B1(_02927_),
    .VDD(VPWR),
    .Y(_01330_),
    .VSS(VGND),
    .A1(net1815),
    .A2(_02926_));
 sg13g2_inv_1 _08722_ (.VDD(VPWR),
    .Y(_02928_),
    .A(\acc_sum.add_renorm0.exp[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08723_ (.Y(_02929_),
    .A(net1819),
    .B(\acc_sum.seg_reg0.q[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08724_ (.B1(_02929_),
    .VDD(VPWR),
    .Y(_01329_),
    .VSS(VGND),
    .A1(net1815),
    .A2(_02928_));
 sg13g2_inv_1 _08725_ (.VDD(VPWR),
    .Y(_02930_),
    .A(\acc_sum.add_renorm0.exp[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08726_ (.Y(_02931_),
    .A(net1815),
    .B(\acc_sum.seg_reg0.q[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08727_ (.B1(_02931_),
    .VDD(VPWR),
    .Y(_01328_),
    .VSS(VGND),
    .A1(net1815),
    .A2(_02930_));
 sg13g2_inv_1 _08728_ (.VDD(VPWR),
    .Y(_02932_),
    .A(\acc_sum.add_renorm0.exp[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08729_ (.Y(_02933_),
    .A(net1815),
    .B(\acc_sum.seg_reg0.q[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08730_ (.B1(_02933_),
    .VDD(VPWR),
    .Y(_01327_),
    .VSS(VGND),
    .A1(net1815),
    .A2(_02932_));
 sg13g2_nor2_1 _08731_ (.A(\acc_sum.exp_mant_logic0.a[15] ),
    .B(\acc_sum.reg1en.d[0] ),
    .Y(_02934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08732_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01723_),
    .A2(\acc_sum.reg1en.d[0] ),
    .Y(_01326_),
    .B1(_02934_));
 sg13g2_inv_1 _08733_ (.VDD(VPWR),
    .Y(_02935_),
    .A(\acc_sum.exp_mant_logic0.a[14] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08734_ (.Y(_02936_),
    .A(\acc[14] ),
    .B(net1901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08735_ (.B1(_02936_),
    .VDD(VPWR),
    .Y(_01325_),
    .VSS(VGND),
    .A1(net1903),
    .A2(_02935_));
 sg13g2_inv_2 _08736_ (.Y(_02937_),
    .A(\acc_sum.exp_mant_logic0.a[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08737_ (.Y(_02938_),
    .A(\acc[13] ),
    .B(net1901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08738_ (.B1(_02938_),
    .VDD(VPWR),
    .Y(_01324_),
    .VSS(VGND),
    .A1(net1904),
    .A2(_02937_));
 sg13g2_inv_1 _08739_ (.VDD(VPWR),
    .Y(_02939_),
    .A(\acc_sum.exp_mant_logic0.a[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08740_ (.Y(_02940_),
    .A(\acc[12] ),
    .B(net1901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08741_ (.B1(_02940_),
    .VDD(VPWR),
    .Y(_01323_),
    .VSS(VGND),
    .A1(net1904),
    .A2(_02939_));
 sg13g2_inv_1 _08742_ (.VDD(VPWR),
    .Y(_02941_),
    .A(\acc_sum.exp_mant_logic0.a[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08743_ (.Y(_02942_),
    .A(\acc[11] ),
    .B(net1901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08744_ (.B1(_02942_),
    .VDD(VPWR),
    .Y(_01322_),
    .VSS(VGND),
    .A1(net1903),
    .A2(_02941_));
 sg13g2_inv_1 _08745_ (.VDD(VPWR),
    .Y(_02943_),
    .A(\acc_sum.exp_mant_logic0.a[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08746_ (.Y(_02944_),
    .A(\acc[10] ),
    .B(net1898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08747_ (.B1(_02944_),
    .VDD(VPWR),
    .Y(_01321_),
    .VSS(VGND),
    .A1(net1900),
    .A2(_02943_));
 sg13g2_inv_1 _08748_ (.VDD(VPWR),
    .Y(_02945_),
    .A(\acc_sum.exp_mant_logic0.a[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08749_ (.Y(_02946_),
    .A(\acc[9] ),
    .B(net1897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08750_ (.B1(_02946_),
    .VDD(VPWR),
    .Y(_01320_),
    .VSS(VGND),
    .A1(net1898),
    .A2(_02945_));
 sg13g2_inv_1 _08751_ (.VDD(VPWR),
    .Y(_02947_),
    .A(\acc_sum.exp_mant_logic0.a[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08752_ (.Y(_02948_),
    .A(\acc[8] ),
    .B(net1900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08753_ (.B1(_02948_),
    .VDD(VPWR),
    .Y(_01319_),
    .VSS(VGND),
    .A1(net1900),
    .A2(_02947_));
 sg13g2_inv_2 _08754_ (.Y(_02949_),
    .A(\acc_sum.exp_mant_logic0.a[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08755_ (.Y(_02950_),
    .A(\acc[7] ),
    .B(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08756_ (.B1(_02950_),
    .VDD(VPWR),
    .Y(_01318_),
    .VSS(VGND),
    .A1(net1898),
    .A2(_02949_));
 sg13g2_inv_2 _08757_ (.Y(_02951_),
    .A(\acc_sum.exp_mant_logic0.a[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08758_ (.Y(_02952_),
    .A(\acc[6] ),
    .B(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08759_ (.B1(_02952_),
    .VDD(VPWR),
    .Y(_01317_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_02951_));
 sg13g2_inv_2 _08760_ (.Y(_02953_),
    .A(\acc_sum.exp_mant_logic0.a[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08761_ (.Y(_02954_),
    .A(\acc[5] ),
    .B(net1901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08762_ (.B1(_02954_),
    .VDD(VPWR),
    .Y(_01316_),
    .VSS(VGND),
    .A1(net1905),
    .A2(_02953_));
 sg13g2_inv_1 _08763_ (.VDD(VPWR),
    .Y(_02955_),
    .A(\acc_sum.exp_mant_logic0.a[4] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08764_ (.Y(_02956_),
    .A(\acc[4] ),
    .B(net1897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08765_ (.B1(_02956_),
    .VDD(VPWR),
    .Y(_01315_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_02955_));
 sg13g2_inv_2 _08766_ (.Y(_02957_),
    .A(\acc_sum.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08767_ (.Y(_02958_),
    .A(\acc[3] ),
    .B(net1897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08768_ (.B1(_02958_),
    .VDD(VPWR),
    .Y(_01314_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_02957_));
 sg13g2_inv_2 _08769_ (.Y(_02959_),
    .A(\acc_sum.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08770_ (.Y(_02960_),
    .A(\acc[2] ),
    .B(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08771_ (.B1(_02960_),
    .VDD(VPWR),
    .Y(_01313_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_02959_));
 sg13g2_inv_1 _08772_ (.VDD(VPWR),
    .Y(_02961_),
    .A(\acc_sum.exp_mant_logic0.a[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08773_ (.Y(_02962_),
    .A(\acc[1] ),
    .B(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08774_ (.B1(_02962_),
    .VDD(VPWR),
    .Y(_01312_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_02961_));
 sg13g2_inv_2 _08775_ (.Y(_02963_),
    .A(\acc_sum.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08776_ (.Y(_02964_),
    .A(\acc[0] ),
    .B(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08777_ (.B1(_02964_),
    .VDD(VPWR),
    .Y(_01311_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_02963_));
 sg13g2_inv_1 _08778_ (.VDD(VPWR),
    .Y(_02965_),
    .A(\acc_sub.reg3en.q[0] ),
    .VSS(VGND));
 sg13g2_nand2_2 _08779_ (.Y(_02966_),
    .A(\acc_sub.add_renorm0.mantisa[3] ),
    .B(\acc_sub.add_renorm0.mantisa[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08780_ (.Y(_02967_),
    .A(\acc_sub.add_renorm0.mantisa[4] ),
    .B(_02966_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1756 (.A(_05573_),
    .X(net1756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08782_ (.VDD(VPWR),
    .Y(_02969_),
    .A(_02966_),
    .VSS(VGND));
 sg13g2_nand3_1 _08783_ (.B(\acc_sub.add_renorm0.mantisa[5] ),
    .C(\acc_sub.add_renorm0.mantisa[4] ),
    .A(_02969_),
    .Y(_02970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08784_ (.Y(_02971_),
    .A(\acc_sub.add_renorm0.mantisa[6] ),
    .B(_02970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout93 (.A(net141),
    .X(net93),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08786_ (.VDD(VPWR),
    .Y(_02973_),
    .A(_02971_),
    .VSS(VGND));
 sg13g2_inv_1 _08787_ (.VDD(VPWR),
    .Y(_02974_),
    .A(\acc_sub.add_renorm0.mantisa[9] ),
    .VSS(VGND));
 sg13g2_inv_1 _08788_ (.VDD(VPWR),
    .Y(_02975_),
    .A(\acc_sub.add_renorm0.mantisa[6] ),
    .VSS(VGND));
 sg13g2_nor2_1 _08789_ (.A(_02975_),
    .B(_02970_),
    .Y(_02976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08790_ (.B(\acc_sub.add_renorm0.mantisa[8] ),
    .C(\acc_sub.add_renorm0.mantisa[7] ),
    .A(_02976_),
    .Y(_02977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08791_ (.A(_02974_),
    .B(_02977_),
    .Y(_02978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08792_ (.A(\acc_sub.add_renorm0.mantisa[10] ),
    .B(_02978_),
    .Y(_02979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1724 (.A(_07027_),
    .X(net1724),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08794_ (.Y(_02981_),
    .A(_02977_),
    .B(_02974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08795_ (.Y(_02982_),
    .A(\acc_sub.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08796_ (.B(\acc_sub.add_renorm0.mantisa[5] ),
    .C(\acc_sub.add_renorm0.mantisa[4] ),
    .A(\acc_sub.add_renorm0.mantisa[6] ),
    .Y(_02983_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\acc_sub.add_renorm0.mantisa[3] ));
 sg13g2_nor3_1 _08797_ (.A(_01647_),
    .B(_02982_),
    .C(_02983_),
    .Y(_02984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08798_ (.VDD(VPWR),
    .Y(_02985_),
    .A(\acc_sub.add_renorm0.mantisa[2] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _08799_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_01700_),
    .A2(_01707_),
    .Y(_02986_),
    .B1(_02985_));
 sg13g2_nor2_1 _08800_ (.A(_02969_),
    .B(_02986_),
    .Y(_02987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08801_ (.VDD(VPWR),
    .Y(_02988_),
    .A(_02987_),
    .VSS(VGND));
 sg13g2_nand3_1 _08802_ (.B(\acc_sub.add_renorm0.mantisa[9] ),
    .C(_02988_),
    .A(_02984_),
    .Y(_02989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08803_ (.Y(_02990_),
    .A(_02981_),
    .B(_02989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08804_ (.Y(_02991_),
    .A(net1704),
    .B(_02990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08805_ (.Y(_02992_),
    .A(_02976_),
    .B(\acc_sub.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08806_ (.Y(_02993_),
    .A(_02992_),
    .B(_01647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _08807_ (.A(_02993_),
    .B(_02977_),
    .X(_02994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08808_ (.Y(_02995_),
    .A(_02994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08809_ (.Y(_02996_),
    .A(_02982_),
    .B(_02976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08810_ (.Y(_02997_),
    .A(_02996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08811_ (.Y(_02998_),
    .A(_02995_),
    .B(_02997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _08812_ (.A(_02973_),
    .B(_02991_),
    .C(_02998_),
    .Y(_02999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08813_ (.B1(_02966_),
    .VDD(VPWR),
    .Y(_03000_),
    .VSS(VGND),
    .A1(\acc_sub.add_renorm0.mantisa[3] ),
    .A2(_02986_));
 sg13g2_inv_4 _08814_ (.A(_03000_),
    .Y(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08815_ (.Y(_03002_),
    .A(\acc_sub.add_renorm0.mantisa[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08816_ (.A(_02966_),
    .B_N(\acc_sub.add_renorm0.mantisa[4] ),
    .Y(_03003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08817_ (.Y(_03004_),
    .A(_03002_),
    .B(_03003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1763 (.A(_03988_),
    .X(net1763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08819_ (.VDD(VPWR),
    .Y(_03006_),
    .A(_03004_),
    .VSS(VGND));
 sg13g2_nor4_1 _08820_ (.A(_02971_),
    .B(_03006_),
    .C(_02991_),
    .D(_02998_),
    .Y(_03007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08821_ (.Y(_03008_),
    .B1(_03001_),
    .B2(_03007_),
    .A2(_02999_),
    .A1(_02967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _08822_ (.A(net1704),
    .Y(_03009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08823_ (.A(_02990_),
    .B(_03009_),
    .Y(_03010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08824_ (.A(_02979_),
    .B(_02995_),
    .Y(_03011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03010_),
    .A2(_02996_),
    .Y(_03012_),
    .B1(_03011_));
 sg13g2_inv_2 _08826_ (.Y(_03013_),
    .A(_02990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _08827_ (.A(_02995_),
    .B(_03013_),
    .C(_03009_),
    .Y(_03014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08829_ (.B(net1704),
    .C(_02990_),
    .A(_02995_),
    .Y(_03016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08830_ (.A(_02997_),
    .B(_03016_),
    .Y(_03017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08831_ (.Y(_03018_),
    .B1(_03004_),
    .B2(_03017_),
    .A2(_02971_),
    .A1(_03014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08832_ (.B(_03012_),
    .C(_03018_),
    .A(_03008_),
    .Y(_03019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08833_ (.Y(_03020_),
    .A(net1788),
    .B(\acc_sub.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08834_ (.B1(_03020_),
    .VDD(VPWR),
    .Y(_03021_),
    .VSS(VGND),
    .A1(net1788),
    .A2(_01647_));
 sg13g2_nand2_1 _08835_ (.Y(_03022_),
    .A(_03002_),
    .B(net1789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08836_ (.B1(_03022_),
    .VDD(VPWR),
    .Y(_03023_),
    .VSS(VGND),
    .A1(net1789),
    .A2(\acc_sub.add_renorm0.mantisa[4] ));
 sg13g2_inv_1 _08837_ (.VDD(VPWR),
    .Y(_03024_),
    .A(net1788),
    .VSS(VGND));
 sg13g2_inv_1 _08838_ (.VDD(VPWR),
    .Y(_03025_),
    .A(\acc_sub.add_renorm0.mantisa[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _08839_ (.Y(_03026_),
    .A(_03024_),
    .B(_03025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08840_ (.B1(_03026_),
    .VDD(VPWR),
    .Y(_03027_),
    .VSS(VGND),
    .A1(_03024_),
    .A2(\acc_sub.add_renorm0.mantisa[4] ));
 sg13g2_buf_2 place1745 (.A(_04268_),
    .X(net1745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08842_ (.A(\acc_sub.add_renorm0.mantisa[11] ),
    .B(\acc_sub.add_renorm0.mantisa[2] ),
    .Y(_03029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08843_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1788),
    .A2(_03025_),
    .Y(_03030_),
    .B1(_03029_));
 sg13g2_inv_1 _08844_ (.VDD(VPWR),
    .Y(_03031_),
    .A(_03030_),
    .VSS(VGND));
 sg13g2_nor3_1 _08845_ (.A(_03023_),
    .B(_03027_),
    .C(_03031_),
    .Y(_03032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08846_ (.Y(_03033_),
    .A(net1789),
    .B(\acc_sub.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08847_ (.B1(_03033_),
    .VDD(VPWR),
    .Y(_03034_),
    .VSS(VGND),
    .A1(net1789),
    .A2(_03002_));
 sg13g2_nand2_1 _08848_ (.Y(_03035_),
    .A(_03032_),
    .B(_03034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08849_ (.VDD(VPWR),
    .Y(_03036_),
    .A(_03035_),
    .VSS(VGND));
 sg13g2_nand2_1 _08850_ (.Y(_03037_),
    .A(net1789),
    .B(\acc_sub.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08851_ (.B1(_03037_),
    .VDD(VPWR),
    .Y(_03038_),
    .VSS(VGND),
    .A1(net1789),
    .A2(_02975_));
 sg13g2_buf_2 place1767 (.A(_03983_),
    .X(net1767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08853_ (.Y(_03040_),
    .A(net1789),
    .B(\acc_sub.add_renorm0.mantisa[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08854_ (.B1(_03040_),
    .VDD(VPWR),
    .Y(_03041_),
    .VSS(VGND),
    .A1(net1789),
    .A2(_02982_));
 sg13g2_and3_2 _08855_ (.X(_03042_),
    .A(_03036_),
    .B(_03038_),
    .C(_03041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1708 (.A(_02652_),
    .X(net1708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08857_ (.Y(_03044_),
    .A(_03021_),
    .B(_03042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08858_ (.A(net1787),
    .B(_03044_),
    .Y(_03045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08859_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03045_),
    .Y(_03046_),
    .A2(net1787),
    .A1(_03019_));
 sg13g2_a21oi_1 _08860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03036_),
    .A2(_03038_),
    .Y(_03047_),
    .B1(_03041_));
 sg13g2_nor3_1 _08861_ (.A(\acc_sub.seg_reg1.q[21] ),
    .B(_03047_),
    .C(_03042_),
    .Y(_03048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08862_ (.Y(_03049_),
    .A(_03010_),
    .B(_02971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08863_ (.B1(_03049_),
    .VDD(VPWR),
    .Y(_03050_),
    .VSS(VGND),
    .A1(_02979_),
    .A2(_02997_));
 sg13g2_a221oi_1 _08864_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_02967_),
    .C1(_03050_),
    .B1(_03017_),
    .A1(_03014_),
    .Y(_03051_),
    .A2(_03004_));
 sg13g2_nand2_1 _08865_ (.Y(_03052_),
    .A(_02999_),
    .B(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03051_),
    .A2(_03052_),
    .Y(_03053_),
    .B1(net1785));
 sg13g2_nor2_2 _08867_ (.A(_03048_),
    .B(_03053_),
    .Y(_03054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08868_ (.A(_01490_),
    .B(_02979_),
    .Y(_03055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08869_ (.Y(_03056_),
    .B1(_03024_),
    .B2(_01707_),
    .A2(\acc_sub.add_renorm0.mantisa[3] ),
    .A1(_02985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08870_ (.A(\acc_sub.add_renorm0.mantisa[1] ),
    .B(_03029_),
    .C(_03056_),
    .Y(_03057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08871_ (.A(_03031_),
    .B(_03057_),
    .Y(_03058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08872_ (.VDD(VPWR),
    .Y(_03059_),
    .A(_03058_),
    .VSS(VGND));
 sg13g2_nor2_1 _08873_ (.A(_03027_),
    .B(_03031_),
    .Y(_03060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08874_ (.A(_03060_),
    .B(_03058_),
    .Y(_03061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08875_ (.A(net1790),
    .B(\acc_sub.add_renorm0.mantisa[10] ),
    .Y(_03062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08876_ (.VDD(VPWR),
    .Y(_03063_),
    .A(_03041_),
    .VSS(VGND));
 sg13g2_nand2_1 _08877_ (.Y(_03064_),
    .A(_03034_),
    .B(_03038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _08878_ (.A(_03023_),
    .B(_03027_),
    .C(_03063_),
    .D(_03064_),
    .Y(_03065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08879_ (.Y(_03066_),
    .A(net1788),
    .B(\acc_sub.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08880_ (.B1(_03066_),
    .VDD(VPWR),
    .Y(_03067_),
    .VSS(VGND),
    .A1(net1788),
    .A2(_02974_));
 sg13g2_nand3_1 _08881_ (.B(_03067_),
    .C(_03021_),
    .A(_03065_),
    .Y(_03068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1749 (.A(net1748),
    .X(net1749),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _08883_ (.A(_03061_),
    .B(_03062_),
    .C(_03068_),
    .Y(_03070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03059_),
    .A2(_03027_),
    .Y(_03071_),
    .B1(_03070_));
 sg13g2_o21ai_1 _08885_ (.B1(_03060_),
    .VDD(VPWR),
    .Y(_03072_),
    .VSS(VGND),
    .A1(_03062_),
    .A2(_03068_));
 sg13g2_and2_1 _08886_ (.A(_03072_),
    .B(_01490_),
    .X(_03073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08887_ (.Y(_03074_),
    .B1(_03071_),
    .B2(_03073_),
    .A2(_03055_),
    .A1(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08888_ (.A(_03062_),
    .B(_03030_),
    .Y(_03075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08889_ (.Y(_03076_),
    .A(_03062_),
    .B(_03068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _08890_ (.A(_03076_),
    .B_N(_03057_),
    .Y(_03077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08891_ (.A(_03059_),
    .B(_03076_),
    .Y(_03078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08892_ (.A(_03075_),
    .B(_03077_),
    .C(_03078_),
    .Y(_03079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08893_ (.VDD(VPWR),
    .Y(_03080_),
    .A(_03070_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03079_),
    .A2(_03080_),
    .Y(_03081_),
    .B1(net1787));
 sg13g2_nor2_1 _08895_ (.A(_03006_),
    .B(_02971_),
    .Y(_03082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08896_ (.Y(_03083_),
    .A(_02973_),
    .B(_03006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08897_ (.A(_03000_),
    .B(_02967_),
    .C(_03083_),
    .Y(_03084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08898_ (.A(_02991_),
    .B(_02998_),
    .Y(_03085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08899_ (.B1(_03085_),
    .VDD(VPWR),
    .Y(_03086_),
    .VSS(VGND),
    .A1(_03082_),
    .A2(_03084_));
 sg13g2_inv_1 _08900_ (.VDD(VPWR),
    .Y(_03087_),
    .A(_03017_),
    .VSS(VGND));
 sg13g2_inv_1 _08901_ (.VDD(VPWR),
    .Y(_03088_),
    .A(_03010_),
    .VSS(VGND));
 sg13g2_nand3_1 _08902_ (.B(_03087_),
    .C(_03088_),
    .A(_03086_),
    .Y(_03089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1704 (.A(_02979_),
    .X(net1704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08904_ (.VDD(VPWR),
    .Y(_03091_),
    .A(_03089_),
    .VSS(VGND));
 sg13g2_inv_1 _08905_ (.VDD(VPWR),
    .Y(_03092_),
    .A(_02967_),
    .VSS(VGND));
 sg13g2_nor3_1 _08906_ (.A(_03092_),
    .B(_02996_),
    .C(_03083_),
    .Y(_03093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _08907_ (.A(_03016_),
    .B_N(_03093_),
    .Y(_03094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_5_4__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08909_ (.A(_03014_),
    .B(_03094_),
    .Y(_03096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08910_ (.Y(_03097_),
    .A(_03096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08911_ (.A(_03013_),
    .B(_02973_),
    .C(_02998_),
    .Y(_03098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08912_ (.A(_03009_),
    .B(_03098_),
    .Y(_03099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08913_ (.VDD(VPWR),
    .Y(_03100_),
    .A(_03099_),
    .VSS(VGND));
 sg13g2_nor2_1 _08914_ (.A(_03097_),
    .B(_03100_),
    .Y(_03101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08915_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03091_),
    .A2(_03101_),
    .Y(_03102_),
    .B1(net1785));
 sg13g2_nor2_1 _08916_ (.A(_03081_),
    .B(_03102_),
    .Y(_03103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08917_ (.B(_03054_),
    .C(_03074_),
    .A(_03046_),
    .Y(_03104_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03103_));
 sg13g2_a22oi_1 _08918_ (.Y(_03105_),
    .B1(_02967_),
    .B2(_03007_),
    .A2(_02999_),
    .A1(_03004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08919_ (.B1(_03013_),
    .VDD(VPWR),
    .Y(_03106_),
    .VSS(VGND),
    .A1(_02994_),
    .A2(_03009_));
 sg13g2_a22oi_1 _08920_ (.Y(_03107_),
    .B1(_02971_),
    .B2(_03017_),
    .A2(_03014_),
    .A1(_02996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08921_ (.Y(_03108_),
    .A(_03094_),
    .B(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _08922_ (.B(_03106_),
    .C(_03107_),
    .A(_03105_),
    .Y(_03109_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03108_));
 sg13g2_nand2_1 _08923_ (.Y(_03110_),
    .A(_03042_),
    .B(_03021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _08924_ (.B(_03110_),
    .A(_03067_),
    .X(_03111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08925_ (.A(\acc_sub.seg_reg1.q[21] ),
    .B(_03111_),
    .Y(_03112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _08926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03109_),
    .A2(net1787),
    .Y(_03113_),
    .B1(_03112_));
 sg13g2_xnor2_1 _08927_ (.Y(_03114_),
    .A(_03038_),
    .B(_03035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _08928_ (.Y(_03115_),
    .B1(_03004_),
    .B2(_03010_),
    .A2(_02971_),
    .A1(_03009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08929_ (.Y(_03116_),
    .A(_03017_),
    .B(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08930_ (.Y(_03117_),
    .A(_03014_),
    .B(_02967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08931_ (.B(_03116_),
    .C(_03117_),
    .A(_03115_),
    .Y(_03118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _08932_ (.A0(_03114_),
    .A1(_03118_),
    .S(\acc_sub.seg_reg1.q[21] ),
    .X(_03119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08933_ (.Y(_03120_),
    .A(_03119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08934_ (.Y(_03121_),
    .A(_03010_),
    .B(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08935_ (.B1(_03121_),
    .VDD(VPWR),
    .Y(_03122_),
    .VSS(VGND),
    .A1(_02979_),
    .A2(_03092_));
 sg13g2_nor2b_1 _08936_ (.A(_03060_),
    .B_N(_03023_),
    .Y(_03123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08937_ (.A(\acc_sub.seg_reg1.q[21] ),
    .B(_03032_),
    .C(_03123_),
    .Y(_03124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08938_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03124_),
    .Y(_03125_),
    .A2(net1787),
    .A1(_03122_));
 sg13g2_nand2_1 _08939_ (.Y(_03126_),
    .A(_03014_),
    .B(_03001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08940_ (.Y(_03127_),
    .A(_03009_),
    .B(_03004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08941_ (.Y(_03128_),
    .A(_03010_),
    .B(_02967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _08942_ (.B(_03127_),
    .C(_03128_),
    .A(_03126_),
    .Y(_03129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08943_ (.A(_03034_),
    .B(_03032_),
    .Y(_03130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _08944_ (.A(\acc_sub.seg_reg1.q[21] ),
    .B(_03130_),
    .C(_03036_),
    .Y(_03131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08945_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03131_),
    .Y(_03132_),
    .A2(\acc_sub.seg_reg1.q[21] ),
    .A1(_03129_));
 sg13g2_nand4_1 _08946_ (.B(_03120_),
    .C(_03125_),
    .A(_03113_),
    .Y(_03133_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03132_));
 sg13g2_nor2_1 _08947_ (.A(_03104_),
    .B(_03133_),
    .Y(_03134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _08948_ (.A(_02965_),
    .B(_03134_),
    .Y(_03135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08949_ (.Y(_03136_),
    .A(_03135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08950_ (.Y(_03137_),
    .A(net1773),
    .B(\acc_sub.y[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _08951_ (.B1(_03137_),
    .VDD(VPWR),
    .Y(_01310_),
    .VSS(VGND),
    .A1(_01498_),
    .A2(_03136_));
 sg13g2_inv_1 _08952_ (.VDD(VPWR),
    .Y(_03138_),
    .A(\acc_sub.y[14] ),
    .VSS(VGND));
 sg13g2_nand3_1 _08953_ (.B(\acc_sub.add_renorm0.exp[1] ),
    .C(\acc_sub.add_renorm0.exp[0] ),
    .A(\acc_sub.add_renorm0.exp[2] ),
    .Y(_03139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08954_ (.A(_01717_),
    .B(_03139_),
    .Y(_03140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08955_ (.Y(_03141_),
    .A(_03140_),
    .B(\acc_sub.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08956_ (.A(_01713_),
    .B(_03141_),
    .Y(_03142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08957_ (.Y(_03143_),
    .A(_03142_),
    .B(\acc_sub.add_renorm0.exp[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08958_ (.Y(_03144_),
    .A(_01709_),
    .B(_03143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _08959_ (.Y(_03145_),
    .A(_02978_),
    .B(\acc_sub.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _08960_ (.Y(_03146_),
    .A(_03145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout129 (.A(net140),
    .X(net129),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08962_ (.A(\acc_sub.add_renorm0.exp[7] ),
    .B(net1699),
    .Y(_03148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08963_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03148_),
    .Y(_03149_),
    .A2(net1699),
    .A1(_03144_));
 sg13g2_xnor2_1 _08964_ (.Y(_03150_),
    .A(_01711_),
    .B(_03142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08965_ (.VDD(VPWR),
    .Y(_03151_),
    .A(_03150_),
    .VSS(VGND));
 sg13g2_nor2_1 _08966_ (.A(\acc_sub.add_renorm0.exp[6] ),
    .B(net1699),
    .Y(_03152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08967_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03152_),
    .Y(_03153_),
    .A2(_03151_),
    .A1(net1699));
 sg13g2_xnor2_1 _08968_ (.Y(_03154_),
    .A(\acc_sub.add_renorm0.exp[3] ),
    .B(_03139_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08969_ (.VDD(VPWR),
    .Y(_03155_),
    .A(_03154_),
    .VSS(VGND));
 sg13g2_nor2_1 _08970_ (.A(\acc_sub.add_renorm0.exp[3] ),
    .B(net1699),
    .Y(_03156_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08971_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03156_),
    .Y(_03157_),
    .A2(_03155_),
    .A1(net1699));
 sg13g2_nand2_1 _08972_ (.Y(_03158_),
    .A(_03085_),
    .B(_03084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08973_ (.Y(_03159_),
    .A(_03146_),
    .B(\acc_sub.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08974_ (.Y(_03160_),
    .A(_01721_),
    .B(_03159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08975_ (.VDD(VPWR),
    .Y(_03161_),
    .A(_03160_),
    .VSS(VGND));
 sg13g2_a21oi_1 _08976_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03087_),
    .A2(_03158_),
    .Y(_03162_),
    .B1(_03161_));
 sg13g2_nand3_1 _08977_ (.B(_03087_),
    .C(_03158_),
    .A(_03161_),
    .Y(_03163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08978_ (.Y(_03164_),
    .B(_03163_),
    .A_N(_03162_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08979_ (.Y(_03165_),
    .A(\acc_sub.add_renorm0.exp[0] ),
    .B(_03145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _08980_ (.Y(_03166_),
    .B(_03165_),
    .A_N(_03164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08981_ (.Y(_03167_),
    .A(_03166_),
    .B(_03163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08982_ (.VDD(VPWR),
    .Y(_03168_),
    .A(\acc_sub.add_renorm0.exp[0] ),
    .VSS(VGND));
 sg13g2_o21ai_1 _08983_ (.B1(_01719_),
    .VDD(VPWR),
    .Y(_03169_),
    .VSS(VGND),
    .A1(_01721_),
    .A2(_03168_));
 sg13g2_and2_1 _08984_ (.A(_03169_),
    .B(_03139_),
    .X(_03170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08985_ (.VDD(VPWR),
    .Y(_03171_),
    .A(_03170_),
    .VSS(VGND));
 sg13g2_nor2_1 _08986_ (.A(\acc_sub.add_renorm0.exp[2] ),
    .B(_03146_),
    .Y(_03172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08987_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03172_),
    .Y(_03173_),
    .A2(_03171_),
    .A1(_03146_));
 sg13g2_buf_1 place1715 (.A(_06907_),
    .X(net1715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08989_ (.VDD(VPWR),
    .Y(_03175_),
    .A(_03173_),
    .VSS(VGND));
 sg13g2_xnor2_1 _08990_ (.Y(_03176_),
    .A(_03175_),
    .B(_03086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08991_ (.Y(_03177_),
    .A(_03167_),
    .B(_03176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08992_ (.Y(_03178_),
    .A(_03086_),
    .B(_03173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _08993_ (.Y(_03179_),
    .A(_03177_),
    .B(_03178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08994_ (.A(_03157_),
    .B(_03179_),
    .Y(_03180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _08995_ (.Y(_03181_),
    .A(\acc_sub.add_renorm0.exp[5] ),
    .B(_03141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _08996_ (.A(_03181_),
    .B(_03145_),
    .Y(_03182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _08997_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03182_),
    .Y(_03183_),
    .A2(_03145_),
    .A1(_01713_));
 sg13g2_xnor2_1 _08998_ (.Y(_03184_),
    .A(_01715_),
    .B(_03140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _08999_ (.VDD(VPWR),
    .Y(_03185_),
    .A(_03184_),
    .VSS(VGND));
 sg13g2_nor2_1 _09000_ (.A(\acc_sub.add_renorm0.exp[4] ),
    .B(net1699),
    .Y(_03186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09001_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03186_),
    .Y(_03187_),
    .A2(_03185_),
    .A1(net1699));
 sg13g2_nor2_1 _09002_ (.A(_03183_),
    .B(_03187_),
    .Y(_03188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09003_ (.Y(_03189_),
    .A(_03180_),
    .B(_03188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09004_ (.A(_03153_),
    .B(_03189_),
    .Y(_03190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09005_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03190_),
    .A2(_03149_),
    .Y(_03191_),
    .B1(_03091_));
 sg13g2_o21ai_1 _09006_ (.B1(_03191_),
    .VDD(VPWR),
    .Y(_03192_),
    .VSS(VGND),
    .A1(_03149_),
    .A2(_03190_));
 sg13g2_inv_1 _09007_ (.VDD(VPWR),
    .Y(_03193_),
    .A(_03149_),
    .VSS(VGND));
 sg13g2_nor3_1 _09008_ (.A(_03009_),
    .B(_03157_),
    .C(_03173_),
    .Y(_03194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09009_ (.VDD(VPWR),
    .Y(_03195_),
    .A(_03187_),
    .VSS(VGND));
 sg13g2_nand2_1 _09010_ (.Y(_03196_),
    .A(_03194_),
    .B(_03195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09011_ (.A(_03183_),
    .B(_03196_),
    .Y(_03197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09012_ (.VDD(VPWR),
    .Y(_03198_),
    .A(_03153_),
    .VSS(VGND));
 sg13g2_nand2_1 _09013_ (.Y(_03199_),
    .A(_03197_),
    .B(_03198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09014_ (.Y(_03200_),
    .A(_03193_),
    .B(_03199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09015_ (.A(_03099_),
    .B(_03200_),
    .Y(_03201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09016_ (.VDD(VPWR),
    .Y(_03202_),
    .A(_03094_),
    .VSS(VGND));
 sg13g2_xor2_1 _09017_ (.B(_03173_),
    .A(_03094_),
    .X(_03203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09018_ (.A(_03160_),
    .B(_03203_),
    .Y(_03204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09019_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03202_),
    .A2(_03173_),
    .Y(_03205_),
    .B1(_03204_));
 sg13g2_inv_1 _09020_ (.VDD(VPWR),
    .Y(_03206_),
    .A(_03157_),
    .VSS(VGND));
 sg13g2_nand2_1 _09021_ (.Y(_03207_),
    .A(_03205_),
    .B(_03206_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09022_ (.VDD(VPWR),
    .Y(_03208_),
    .A(_03207_),
    .VSS(VGND));
 sg13g2_nand2_1 _09023_ (.Y(_03209_),
    .A(_03208_),
    .B(_03195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09024_ (.A(_03183_),
    .B(_03209_),
    .Y(_03210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09025_ (.Y(_03211_),
    .A(_03210_),
    .B(_03198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09026_ (.B1(_03097_),
    .VDD(VPWR),
    .Y(_03212_),
    .VSS(VGND),
    .A1(_03193_),
    .A2(_03211_));
 sg13g2_a21oi_1 _09027_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03193_),
    .A2(_03211_),
    .Y(_03213_),
    .B1(_03212_));
 sg13g2_nor3_1 _09028_ (.A(net1785),
    .B(_03201_),
    .C(_03213_),
    .Y(_03214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09029_ (.Y(_03215_),
    .A(_03192_),
    .B(_03214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09030_ (.A(net1791),
    .B(\acc_sub.add_renorm0.exp[7] ),
    .Y(_03216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09031_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03144_),
    .A2(net1791),
    .Y(_03217_),
    .B1(_03216_));
 sg13g2_nor2_1 _09032_ (.A(net1790),
    .B(_01717_),
    .Y(_03218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _09033_ (.A2(net1790),
    .A1(_03154_),
    .B1(_03218_),
    .X(_03219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09034_ (.VDD(VPWR),
    .Y(_03220_),
    .A(_03219_),
    .VSS(VGND));
 sg13g2_nor2_1 _09035_ (.A(net1790),
    .B(_01719_),
    .Y(_03221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _09036_ (.A2(net1790),
    .A1(_03170_),
    .B1(_03221_),
    .X(_03222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09037_ (.VDD(VPWR),
    .Y(_03223_),
    .A(_03222_),
    .VSS(VGND));
 sg13g2_nor2_1 _09038_ (.A(net1790),
    .B(\acc_sub.add_renorm0.exp[0] ),
    .Y(_03224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09039_ (.Y(_03225_),
    .A(net1790),
    .B(\acc_sub.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _09040_ (.A(_03224_),
    .B_N(_03225_),
    .Y(_03226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _09041_ (.A(_03080_),
    .B_N(_03226_),
    .Y(_03227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09042_ (.Y(_03228_),
    .A(_03227_),
    .B(\acc_sub.add_renorm0.exp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09043_ (.A(_03223_),
    .B(_03228_),
    .Y(_03229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09044_ (.VDD(VPWR),
    .Y(_03230_),
    .A(_03229_),
    .VSS(VGND));
 sg13g2_nor2_1 _09045_ (.A(_03220_),
    .B(_03230_),
    .Y(_03231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09046_ (.A(net1791),
    .B(_01715_),
    .Y(_03232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _09047_ (.A2(net1791),
    .A1(_03184_),
    .B1(_03232_),
    .X(_03233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _09048_ (.A(_03231_),
    .B(_03233_),
    .X(_03234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09049_ (.Y(_03235_),
    .A(_03181_),
    .B(net1791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09050_ (.B1(_03235_),
    .VDD(VPWR),
    .Y(_03236_),
    .VSS(VGND),
    .A1(net1791),
    .A2(_01713_));
 sg13g2_nand2_1 _09051_ (.Y(_03237_),
    .A(_03234_),
    .B(_03236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09052_ (.A(net1791),
    .B(\acc_sub.add_renorm0.exp[6] ),
    .Y(_03238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09053_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03151_),
    .A2(net1791),
    .Y(_03239_),
    .B1(_03238_));
 sg13g2_nor2b_1 _09054_ (.A(_03237_),
    .B_N(_03239_),
    .Y(_03240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09055_ (.Y(_03241_),
    .A(_03217_),
    .B(_03240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09056_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1786),
    .A2(_03241_),
    .Y(_03242_),
    .B1(_03136_));
 sg13g2_nand2_1 _09057_ (.Y(_03243_),
    .A(_03215_),
    .B(_03242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09058_ (.B1(_03243_),
    .VDD(VPWR),
    .Y(_01309_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03138_));
 sg13g2_inv_2 _09059_ (.Y(_03244_),
    .A(\acc_sub.y[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09060_ (.VDD(VPWR),
    .Y(_03245_),
    .A(_03189_),
    .VSS(VGND));
 sg13g2_nor2_1 _09061_ (.A(_03198_),
    .B(_03245_),
    .Y(_03246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09062_ (.B1(_03089_),
    .VDD(VPWR),
    .Y(_03247_),
    .VSS(VGND),
    .A1(_03190_),
    .A2(_03246_));
 sg13g2_inv_1 _09063_ (.VDD(VPWR),
    .Y(_03248_),
    .A(_03197_),
    .VSS(VGND));
 sg13g2_nand2_1 _09064_ (.Y(_03249_),
    .A(_03248_),
    .B(_03153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09065_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03249_),
    .A2(_03199_),
    .Y(_03250_),
    .B1(_03099_));
 sg13g2_inv_1 _09066_ (.VDD(VPWR),
    .Y(_03251_),
    .A(_03210_),
    .VSS(VGND));
 sg13g2_nand2_1 _09067_ (.Y(_03252_),
    .A(_03251_),
    .B(_03153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09068_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03252_),
    .A2(_03211_),
    .Y(_03253_),
    .B1(_03096_));
 sg13g2_nor3_1 _09069_ (.A(net1785),
    .B(_03250_),
    .C(_03253_),
    .Y(_03254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09070_ (.Y(_03255_),
    .A(_03247_),
    .B(_03254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _09071_ (.B(_03237_),
    .A(_03239_),
    .X(_03256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09072_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1786),
    .A2(_03256_),
    .Y(_03257_),
    .B1(_03136_));
 sg13g2_nand2_1 _09073_ (.Y(_03258_),
    .A(_03255_),
    .B(_03257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09074_ (.B1(_03258_),
    .VDD(VPWR),
    .Y(_01308_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03244_));
 sg13g2_inv_1 _09075_ (.VDD(VPWR),
    .Y(_03259_),
    .A(\acc_sub.y[12] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _09076_ (.Y(_03260_),
    .A(_03236_),
    .B(_03234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09077_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1786),
    .A2(_03260_),
    .Y(_03261_),
    .B1(_03136_));
 sg13g2_nor3_1 _09078_ (.A(_03187_),
    .B(_03157_),
    .C(_03179_),
    .Y(_03262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _09079_ (.A(_03262_),
    .B_N(_03183_),
    .Y(_03263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09080_ (.B1(_03089_),
    .VDD(VPWR),
    .Y(_03264_),
    .VSS(VGND),
    .A1(_03245_),
    .A2(_03263_));
 sg13g2_nand2_1 _09081_ (.Y(_03265_),
    .A(_03196_),
    .B(_03183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09082_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03248_),
    .A2(_03265_),
    .Y(_03266_),
    .B1(_03099_));
 sg13g2_nand2_1 _09083_ (.Y(_03267_),
    .A(_03209_),
    .B(_03183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09084_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03251_),
    .A2(_03267_),
    .Y(_03268_),
    .B1(_03096_));
 sg13g2_nor3_1 _09085_ (.A(net1785),
    .B(_03266_),
    .C(_03268_),
    .Y(_03269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09086_ (.Y(_03270_),
    .A(_03264_),
    .B(_03269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09087_ (.Y(_03271_),
    .A(_03261_),
    .B(_03270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09088_ (.B1(_03271_),
    .VDD(VPWR),
    .Y(_01307_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03259_));
 sg13g2_inv_2 _09089_ (.Y(_03272_),
    .A(\acc_sub.y[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09090_ (.A(_03195_),
    .B(_03180_),
    .Y(_03273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09091_ (.B1(_03089_),
    .VDD(VPWR),
    .Y(_03274_),
    .VSS(VGND),
    .A1(_03262_),
    .A2(_03273_));
 sg13g2_nand2b_1 _09092_ (.Y(_03275_),
    .B(_03187_),
    .A_N(_03194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _09093_ (.A2(_03196_),
    .A1(_03275_),
    .B1(_03099_),
    .X(_03276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09094_ (.Y(_03277_),
    .A(_03207_),
    .B(_03187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _09095_ (.A2(_03277_),
    .A1(_03209_),
    .B1(_03096_),
    .X(_03278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09096_ (.B(_03276_),
    .C(_03278_),
    .A(_03274_),
    .Y(_03279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09097_ (.Y(_03280_),
    .A(_03233_),
    .B(_03231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09098_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1786),
    .A2(_03280_),
    .Y(_03281_),
    .B1(_03136_));
 sg13g2_o21ai_1 _09099_ (.B1(_03281_),
    .VDD(VPWR),
    .Y(_03282_),
    .VSS(VGND),
    .A1(net1786),
    .A2(_03279_));
 sg13g2_o21ai_1 _09100_ (.B1(_03282_),
    .VDD(VPWR),
    .Y(_01306_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03272_));
 sg13g2_inv_2 _09101_ (.Y(_03283_),
    .A(\acc_sub.y[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09102_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03177_),
    .A2(_03178_),
    .Y(_03284_),
    .B1(_03206_));
 sg13g2_o21ai_1 _09103_ (.B1(_03089_),
    .VDD(VPWR),
    .Y(_03285_),
    .VSS(VGND),
    .A1(_03180_),
    .A2(_03284_));
 sg13g2_a21oi_1 _09104_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03175_),
    .A2(net1704),
    .Y(_03286_),
    .B1(_03206_));
 sg13g2_o21ai_1 _09105_ (.B1(_03100_),
    .VDD(VPWR),
    .Y(_03287_),
    .VSS(VGND),
    .A1(_03194_),
    .A2(_03286_));
 sg13g2_nor2_1 _09106_ (.A(_03206_),
    .B(_03205_),
    .Y(_03288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09107_ (.B1(_03097_),
    .VDD(VPWR),
    .Y(_03289_),
    .VSS(VGND),
    .A1(_03288_),
    .A2(_03208_));
 sg13g2_nand4_1 _09108_ (.B(net1787),
    .C(_03287_),
    .A(_03285_),
    .Y(_03290_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03289_));
 sg13g2_nor2_1 _09109_ (.A(_03219_),
    .B(_03229_),
    .Y(_03291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09110_ (.B1(net1786),
    .VDD(VPWR),
    .Y(_03292_),
    .VSS(VGND),
    .A1(_03291_),
    .A2(_03231_));
 sg13g2_nand3_1 _09111_ (.B(_03135_),
    .C(_03292_),
    .A(_03290_),
    .Y(_03293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09112_ (.B1(_03293_),
    .VDD(VPWR),
    .Y(_01305_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03283_));
 sg13g2_inv_2 _09113_ (.Y(_03294_),
    .A(\acc_sub.y[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03167_),
    .A2(_03176_),
    .Y(_03295_),
    .B1(_03091_));
 sg13g2_o21ai_1 _09115_ (.B1(_03295_),
    .VDD(VPWR),
    .Y(_03296_),
    .VSS(VGND),
    .A1(_03167_),
    .A2(_03176_));
 sg13g2_nand2_1 _09116_ (.Y(_03297_),
    .A(_03173_),
    .B(net1704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09117_ (.B1(_03297_),
    .VDD(VPWR),
    .Y(_03298_),
    .VSS(VGND),
    .A1(_03173_),
    .A2(_02999_));
 sg13g2_a21oi_1 _09118_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03203_),
    .A2(_03160_),
    .Y(_03299_),
    .B1(_03096_));
 sg13g2_nand2b_1 _09119_ (.Y(_03300_),
    .B(_03299_),
    .A_N(_03204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _09120_ (.B(net1787),
    .C(_03298_),
    .A(_03296_),
    .Y(_03301_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03300_));
 sg13g2_a21oi_1 _09121_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03227_),
    .A2(\acc_sub.add_renorm0.exp[1] ),
    .Y(_03302_),
    .B1(_03222_));
 sg13g2_o21ai_1 _09122_ (.B1(net1786),
    .VDD(VPWR),
    .Y(_03303_),
    .VSS(VGND),
    .A1(_03229_),
    .A2(_03302_));
 sg13g2_nand3_1 _09123_ (.B(_03301_),
    .C(_03303_),
    .A(_03135_),
    .Y(_03304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09124_ (.B1(_03304_),
    .VDD(VPWR),
    .Y(_01304_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03294_));
 sg13g2_inv_1 _09125_ (.VDD(VPWR),
    .Y(_03305_),
    .A(\acc_sub.y[8] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _09126_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03080_),
    .A2(_03225_),
    .Y(_03306_),
    .B1(_03224_));
 sg13g2_xnor2_1 _09127_ (.Y(_03307_),
    .A(\acc_sub.add_renorm0.exp[1] ),
    .B(_03306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09128_ (.A(_03161_),
    .B(_03096_),
    .Y(_03308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09129_ (.A(_03160_),
    .B(_03099_),
    .Y(_03309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _09130_ (.A(net1785),
    .B(_03308_),
    .C(_03309_),
    .Y(_03310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09131_ (.Y(_03311_),
    .B(_03164_),
    .A_N(_03165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09132_ (.B(_03089_),
    .C(_03311_),
    .A(_03166_),
    .Y(_03312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09133_ (.Y(_03313_),
    .B1(_03310_),
    .B2(_03312_),
    .A2(_03307_),
    .A1(net1786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09134_ (.Y(_03314_),
    .A(_03135_),
    .B(_03313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09135_ (.B1(_03314_),
    .VDD(VPWR),
    .Y(_01303_),
    .VSS(VGND),
    .A1(net1801),
    .A2(_03305_));
 sg13g2_a21oi_1 _09136_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03101_),
    .A2(_03165_),
    .Y(_03315_),
    .B1(net1785));
 sg13g2_o21ai_1 _09137_ (.B1(_03315_),
    .VDD(VPWR),
    .Y(_03316_),
    .VSS(VGND),
    .A1(_03165_),
    .A2(_03089_));
 sg13g2_nor2_1 _09138_ (.A(net1787),
    .B(_03227_),
    .Y(_03317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09139_ (.B1(_03317_),
    .VDD(VPWR),
    .Y(_03318_),
    .VSS(VGND),
    .A1(_03070_),
    .A2(_03226_));
 sg13g2_a21oi_1 _09140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03316_),
    .A2(_03318_),
    .Y(_03319_),
    .B1(_03136_));
 sg13g2_a21o_1 _09141_ (.A2(\acc_sub.y[7] ),
    .A1(net1773),
    .B1(_03319_),
    .X(_01302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09142_ (.Y(_03320_),
    .A(net1773),
    .B(\acc_sub.y[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09143_ (.B1(_03320_),
    .VDD(VPWR),
    .Y(_01301_),
    .VSS(VGND),
    .A1(net1773),
    .A2(_03113_));
 sg13g2_nor2_1 _09144_ (.A(\acc_sub.reg3en.q[0] ),
    .B(\acc_sub.y[5] ),
    .Y(_03321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09145_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03046_),
    .A2(net1801),
    .Y(_01300_),
    .B1(_03321_));
 sg13g2_nor2_1 _09146_ (.A(net1800),
    .B(\acc_sub.y[4] ),
    .Y(_03322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09147_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03054_),
    .A2(net1800),
    .Y(_01299_),
    .B1(_03322_));
 sg13g2_nor2_1 _09148_ (.A(\acc_sub.reg3en.q[0] ),
    .B(\acc_sub.y[3] ),
    .Y(_03323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09149_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03120_),
    .A2(\acc_sub.reg3en.q[0] ),
    .Y(_01298_),
    .B1(_03323_));
 sg13g2_nor2_1 _09150_ (.A(net1800),
    .B(\acc_sub.y[2] ),
    .Y(_03324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09151_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03132_),
    .A2(net1800),
    .Y(_01297_),
    .B1(_03324_));
 sg13g2_nand2_1 _09152_ (.Y(_03325_),
    .A(net1773),
    .B(\acc_sub.y[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09153_ (.B1(_03325_),
    .VDD(VPWR),
    .Y(_01296_),
    .VSS(VGND),
    .A1(net1773),
    .A2(_03125_));
 sg13g2_nand2_1 _09154_ (.Y(_03326_),
    .A(net1773),
    .B(\acc_sub.y[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09155_ (.B1(_03326_),
    .VDD(VPWR),
    .Y(_01295_),
    .VSS(VGND),
    .A1(net1773),
    .A2(_03074_));
 sg13g2_inv_8 _09156_ (.Y(_03327_),
    .A(\acc_sub.x2[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09157_ (.A(net1896),
    .B(\acc_sum.exp_mant_logic0.b[15] ),
    .Y(_03328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09158_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03327_),
    .A2(net1896),
    .Y(_01294_),
    .B1(_03328_));
 sg13g2_inv_2 _09159_ (.Y(_03329_),
    .A(\acc_sum.exp_mant_logic0.b[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09160_ (.Y(_03330_),
    .A(\acc_sub.x2[14] ),
    .B(net1903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09161_ (.B1(_03330_),
    .VDD(VPWR),
    .Y(_01293_),
    .VSS(VGND),
    .A1(net1903),
    .A2(_03329_));
 sg13g2_inv_1 _09162_ (.VDD(VPWR),
    .Y(_03331_),
    .A(\acc_sum.exp_mant_logic0.b[13] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09163_ (.Y(_03332_),
    .A(\acc_sub.x2[13] ),
    .B(net1903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09164_ (.B1(_03332_),
    .VDD(VPWR),
    .Y(_01292_),
    .VSS(VGND),
    .A1(net1905),
    .A2(_03331_));
 sg13g2_inv_2 _09165_ (.Y(_03333_),
    .A(\acc_sum.exp_mant_logic0.b[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09166_ (.Y(_03334_),
    .A(\acc_sub.x2[12] ),
    .B(net1904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09167_ (.B1(_03334_),
    .VDD(VPWR),
    .Y(_01291_),
    .VSS(VGND),
    .A1(net1904),
    .A2(_03333_));
 sg13g2_inv_1 _09168_ (.VDD(VPWR),
    .Y(_03335_),
    .A(\acc_sum.exp_mant_logic0.b[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09169_ (.Y(_03336_),
    .A(\acc_sub.x2[11] ),
    .B(net1904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09170_ (.B1(_03336_),
    .VDD(VPWR),
    .Y(_01290_),
    .VSS(VGND),
    .A1(net1904),
    .A2(_03335_));
 sg13g2_inv_1 _09171_ (.VDD(VPWR),
    .Y(_03337_),
    .A(\acc_sum.exp_mant_logic0.b[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09172_ (.Y(_03338_),
    .A(\acc_sub.x2[10] ),
    .B(net1900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09173_ (.B1(_03338_),
    .VDD(VPWR),
    .Y(_01289_),
    .VSS(VGND),
    .A1(net1901),
    .A2(_03337_));
 sg13g2_inv_2 _09174_ (.Y(_03339_),
    .A(\acc_sum.exp_mant_logic0.b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09175_ (.Y(_03340_),
    .A(\acc_sub.x2[9] ),
    .B(net1897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09176_ (.B1(_03340_),
    .VDD(VPWR),
    .Y(_01288_),
    .VSS(VGND),
    .A1(net1898),
    .A2(_03339_));
 sg13g2_inv_1 _09177_ (.VDD(VPWR),
    .Y(_03341_),
    .A(\acc_sum.exp_mant_logic0.b[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09178_ (.Y(_03342_),
    .A(\acc_sub.x2[8] ),
    .B(net1897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09179_ (.B1(_03342_),
    .VDD(VPWR),
    .Y(_01287_),
    .VSS(VGND),
    .A1(net1899),
    .A2(_03341_));
 sg13g2_inv_2 _09180_ (.Y(_03343_),
    .A(\acc_sum.exp_mant_logic0.b[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09181_ (.Y(_03344_),
    .A(\acc_sub.x2[7] ),
    .B(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09182_ (.B1(_03344_),
    .VDD(VPWR),
    .Y(_01286_),
    .VSS(VGND),
    .A1(net1898),
    .A2(_03343_));
 sg13g2_inv_2 _09183_ (.Y(_03345_),
    .A(\acc_sum.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09184_ (.Y(_03346_),
    .A(\acc_sub.x2[6] ),
    .B(net1905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09185_ (.B1(_03346_),
    .VDD(VPWR),
    .Y(_01285_),
    .VSS(VGND),
    .A1(net1905),
    .A2(_03345_));
 sg13g2_inv_2 _09186_ (.Y(_03347_),
    .A(\acc_sum.exp_mant_logic0.b[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09187_ (.Y(_03348_),
    .A(\acc_sub.x2[5] ),
    .B(net1905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09188_ (.B1(_03348_),
    .VDD(VPWR),
    .Y(_01284_),
    .VSS(VGND),
    .A1(net1902),
    .A2(_03347_));
 sg13g2_inv_2 _09189_ (.Y(_03349_),
    .A(\acc_sum.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09190_ (.Y(_03350_),
    .A(\acc_sub.x2[4] ),
    .B(net1906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09191_ (.B1(_03350_),
    .VDD(VPWR),
    .Y(_01283_),
    .VSS(VGND),
    .A1(net1906),
    .A2(_03349_));
 sg13g2_inv_2 _09192_ (.Y(_03351_),
    .A(\acc_sum.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09193_ (.Y(_03352_),
    .A(\acc_sub.x2[3] ),
    .B(net1906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09194_ (.B1(_03352_),
    .VDD(VPWR),
    .Y(_01282_),
    .VSS(VGND),
    .A1(net1906),
    .A2(_03351_));
 sg13g2_inv_2 _09195_ (.Y(_03353_),
    .A(\acc_sum.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09196_ (.Y(_03354_),
    .A(\acc_sub.x2[2] ),
    .B(net1906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09197_ (.B1(_03354_),
    .VDD(VPWR),
    .Y(_01281_),
    .VSS(VGND),
    .A1(net1906),
    .A2(_03353_));
 sg13g2_inv_2 _09198_ (.Y(_03355_),
    .A(\acc_sum.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09199_ (.Y(_03356_),
    .A(\acc_sub.x2[1] ),
    .B(net1905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09200_ (.B1(_03356_),
    .VDD(VPWR),
    .Y(_01280_),
    .VSS(VGND),
    .A1(net1902),
    .A2(_03355_));
 sg13g2_inv_2 _09201_ (.Y(_03357_),
    .A(\acc_sum.exp_mant_logic0.b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09202_ (.Y(_03358_),
    .A(\acc_sub.x2[0] ),
    .B(net1906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09203_ (.B1(_03358_),
    .VDD(VPWR),
    .Y(_01279_),
    .VSS(VGND),
    .A1(net1906),
    .A2(_03357_));
 sg13g2_inv_1 _09204_ (.VDD(VPWR),
    .Y(_03359_),
    .A(\fp16_res_pipe.seg_reg1.q[21] ),
    .VSS(VGND));
 sg13g2_buf_2 place1793 (.A(\acc_sub.exp_mant_logic0.a[5] ),
    .X(net1793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _09206_ (.A(\fp16_res_pipe.reg2en.q[0] ),
    .Y(_03361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1792 (.A(\acc_sub.exp_mant_logic0.a[6] ),
    .X(net1792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09208_ (.Y(_03363_),
    .A(\fp16_res_pipe.op_sign_logic0.s_a ),
    .B(\fp16_res_pipe.op_sign_logic0.s_b ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09209_ (.Y(_03364_),
    .A(\fp16_res_pipe.op_sign_logic0.add_sub ),
    .B(_03363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09210_ (.A(_03361_),
    .B(_03364_),
    .Y(_03365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout81 (.A(net93),
    .X(net81),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09212_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03359_),
    .A2(_03361_),
    .Y(_01278_),
    .B1(_03365_));
 sg13g2_inv_1 _09213_ (.VDD(VPWR),
    .Y(_03367_),
    .A(\fp16_res_pipe.seg_reg1.q[20] ),
    .VSS(VGND));
 sg13g2_inv_1 _09214_ (.VDD(VPWR),
    .Y(_03368_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09215_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[10] ),
    .B(_03368_),
    .Y(_03369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09216_ (.VDD(VPWR),
    .Y(_03370_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[8] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09217_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[8] ),
    .B(_03370_),
    .Y(_03371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09218_ (.VDD(VPWR),
    .Y(_03372_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[9] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09219_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[9] ),
    .B(_03372_),
    .Y(_03373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09220_ (.VDD(VPWR),
    .Y(_03374_),
    .A(_03373_),
    .VSS(VGND));
 sg13g2_nand2_1 _09221_ (.Y(_03375_),
    .A(_03372_),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _09222_ (.Y(_03376_),
    .A(_03374_),
    .B(_03375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09223_ (.VDD(VPWR),
    .Y(_03377_),
    .A(_03376_),
    .VSS(VGND));
 sg13g2_inv_1 _09224_ (.VDD(VPWR),
    .Y(_03378_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09225_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[7] ),
    .B(_03378_),
    .Y(_03379_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09226_ (.VDD(VPWR),
    .Y(_03380_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09227_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[7] ),
    .B(_03380_),
    .Y(_03381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09228_ (.A(_03379_),
    .B(_03381_),
    .Y(_03382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09229_ (.VDD(VPWR),
    .Y(_03383_),
    .A(_03382_),
    .VSS(VGND));
 sg13g2_inv_1 _09230_ (.VDD(VPWR),
    .Y(_03384_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[6] ),
    .VSS(VGND));
 sg13g2_nor2_2 _09231_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[6] ),
    .B(_03384_),
    .Y(_03385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09232_ (.VDD(VPWR),
    .Y(_03386_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[6] ),
    .VSS(VGND));
 sg13g2_nor2_2 _09233_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[6] ),
    .B(_03386_),
    .Y(_03387_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09234_ (.A(_03385_),
    .B(_03387_),
    .Y(_03388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09235_ (.VDD(VPWR),
    .Y(_03389_),
    .A(_03388_),
    .VSS(VGND));
 sg13g2_nor2_1 _09236_ (.A(_03383_),
    .B(_03389_),
    .Y(_03390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09237_ (.VDD(VPWR),
    .Y(_03391_),
    .A(_03390_),
    .VSS(VGND));
 sg13g2_inv_1 _09238_ (.VDD(VPWR),
    .Y(_03392_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09239_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[5] ),
    .B(_03392_),
    .Y(_03393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09240_ (.VDD(VPWR),
    .Y(_03394_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09241_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[5] ),
    .B(_03394_),
    .Y(_03395_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09242_ (.A(_03393_),
    .B(_03395_),
    .Y(_03396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09243_ (.Y(_03397_),
    .A(_03396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09244_ (.VDD(VPWR),
    .Y(_03398_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09245_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[3] ),
    .B(_03398_),
    .Y(_03399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09246_ (.VDD(VPWR),
    .Y(_03400_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09247_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[3] ),
    .B(_03400_),
    .Y(_03401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09248_ (.A(_03399_),
    .B(_03401_),
    .Y(_03402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09249_ (.VDD(VPWR),
    .Y(_03403_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09250_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[2] ),
    .B(_03403_),
    .Y(_03404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09251_ (.VDD(VPWR),
    .Y(_03405_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[2] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09252_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[2] ),
    .B(_03405_),
    .Y(_03406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09253_ (.A(_03404_),
    .B(_03406_),
    .Y(_03407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09254_ (.Y(_03408_),
    .A(_03402_),
    .B(_03407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09255_ (.VDD(VPWR),
    .Y(_03409_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[0] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09256_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[0] ),
    .B(_03409_),
    .Y(_03410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09257_ (.VDD(VPWR),
    .Y(_03411_),
    .A(_03410_),
    .VSS(VGND));
 sg13g2_inv_1 _09258_ (.VDD(VPWR),
    .Y(_03412_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09259_ (.Y(_03413_),
    .A(_03412_),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09260_ (.VDD(VPWR),
    .Y(_03414_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09261_ (.Y(_03415_),
    .A(_03414_),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09262_ (.VDD(VPWR),
    .Y(_03416_),
    .A(_03415_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09263_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03411_),
    .A2(_03413_),
    .Y(_03417_),
    .B1(_03416_));
 sg13g2_inv_1 _09264_ (.VDD(VPWR),
    .Y(_03418_),
    .A(_03399_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09265_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03418_),
    .A2(_03406_),
    .Y(_03419_),
    .B1(_03401_));
 sg13g2_o21ai_1 _09266_ (.B1(_03419_),
    .VDD(VPWR),
    .Y(_03420_),
    .VSS(VGND),
    .A1(_03408_),
    .A2(_03417_));
 sg13g2_inv_1 _09267_ (.VDD(VPWR),
    .Y(_03421_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[4] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09268_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[4] ),
    .B(_03421_),
    .Y(_03422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09269_ (.VDD(VPWR),
    .Y(_03423_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[4] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09270_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[4] ),
    .B(_03423_),
    .Y(_03424_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09271_ (.A(_03422_),
    .B(_03424_),
    .Y(_03425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1761 (.A(net1759),
    .X(net1761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09273_ (.Y(_03427_),
    .A(_03420_),
    .B(_03425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09274_ (.VDD(VPWR),
    .Y(_03428_),
    .A(_03393_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09275_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03428_),
    .A2(_03424_),
    .Y(_03429_),
    .B1(_03395_));
 sg13g2_o21ai_1 _09276_ (.B1(_03429_),
    .VDD(VPWR),
    .Y(_03430_),
    .VSS(VGND),
    .A1(_03397_),
    .A2(_03427_));
 sg13g2_inv_1 _09277_ (.VDD(VPWR),
    .Y(_03431_),
    .A(_03430_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09278_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03382_),
    .A2(_03385_),
    .Y(_03432_),
    .B1(_03379_));
 sg13g2_o21ai_1 _09279_ (.B1(_03432_),
    .VDD(VPWR),
    .Y(_03433_),
    .VSS(VGND),
    .A1(_03391_),
    .A2(_03431_));
 sg13g2_inv_1 _09280_ (.VDD(VPWR),
    .Y(_03434_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_b[8] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09281_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_a[8] ),
    .B(_03434_),
    .Y(_03435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09282_ (.A(_03371_),
    .B(_03435_),
    .Y(_03436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09283_ (.VDD(VPWR),
    .Y(_03437_),
    .A(_03436_),
    .VSS(VGND));
 sg13g2_nor2_1 _09284_ (.A(_03376_),
    .B(_03437_),
    .Y(_03438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _09285_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_03438_),
    .C1(_03373_),
    .B1(_03433_),
    .A1(_03371_),
    .Y(_03439_),
    .A2(_03377_));
 sg13g2_nor2_1 _09286_ (.A(_03369_),
    .B(_03439_),
    .Y(_03440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09287_ (.VDD(VPWR),
    .Y(_03441_),
    .A(_03425_),
    .VSS(VGND));
 sg13g2_nor3_1 _09288_ (.A(_03397_),
    .B(_03441_),
    .C(_03408_),
    .Y(_03442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _09289_ (.Y(_03443_),
    .A(_03415_),
    .B(_03413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09290_ (.VDD(VPWR),
    .Y(_03444_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09291_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[10] ),
    .B(_03444_),
    .Y(_03445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09292_ (.A(_03445_),
    .B(_03369_),
    .Y(_03446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09293_ (.VDD(VPWR),
    .Y(_03447_),
    .A(_03446_),
    .VSS(VGND));
 sg13g2_nor2b_1 _09294_ (.A(\fp16_res_pipe.op_sign_logic0.mantisa_b[0] ),
    .B_N(\fp16_res_pipe.op_sign_logic0.mantisa_a[0] ),
    .Y(_03448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09295_ (.VDD(VPWR),
    .Y(_03449_),
    .A(_03448_),
    .VSS(VGND));
 sg13g2_nand2_1 _09296_ (.Y(_03450_),
    .A(_03449_),
    .B(_03411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _09297_ (.A(_03443_),
    .B(_03447_),
    .C(_03450_),
    .Y(_03451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _09298_ (.B(_03451_),
    .C(_03438_),
    .A(_03442_),
    .Y(_03452_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03390_));
 sg13g2_a21oi_2 _09299_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03445_),
    .Y(_03453_),
    .A2(_03452_),
    .A1(_03440_));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1683 (.A(_04052_),
    .X(net1683),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09302_ (.Y(_03456_),
    .A(\fp16_res_pipe.op_sign_logic0.s_b ),
    .B(\fp16_res_pipe.op_sign_logic0.add_sub ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09303_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03453_),
    .A2(_03456_),
    .Y(_03457_),
    .B1(_03361_));
 sg13g2_o21ai_1 _09304_ (.B1(_03457_),
    .VDD(VPWR),
    .Y(_03458_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.op_sign_logic0.s_a ),
    .A2(_03453_));
 sg13g2_o21ai_1 _09305_ (.B1(_03458_),
    .VDD(VPWR),
    .Y(_01277_),
    .VSS(VGND),
    .A1(net1833),
    .A2(_03367_));
 sg13g2_nand2_1 _09306_ (.Y(_03459_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[0] ),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09307_ (.Y(_03460_),
    .B(_03443_),
    .A_N(_03459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09308_ (.B1(_03460_),
    .VDD(VPWR),
    .Y(_03461_),
    .VSS(VGND),
    .A1(_03412_),
    .A2(_03414_));
 sg13g2_nand2b_1 _09309_ (.Y(_03462_),
    .B(_03461_),
    .A_N(_03407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09310_ (.B1(_03462_),
    .VDD(VPWR),
    .Y(_03463_),
    .VSS(VGND),
    .A1(_03405_),
    .A2(_03403_));
 sg13g2_inv_1 _09311_ (.VDD(VPWR),
    .Y(_03464_),
    .A(_03402_),
    .VSS(VGND));
 sg13g2_nand2_1 _09312_ (.Y(_03465_),
    .A(_03463_),
    .B(_03464_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09313_ (.B1(_03465_),
    .VDD(VPWR),
    .Y(_03466_),
    .VSS(VGND),
    .A1(_03400_),
    .A2(_03398_));
 sg13g2_nand2_1 _09314_ (.Y(_03467_),
    .A(_03466_),
    .B(_03441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09315_ (.B1(_03467_),
    .VDD(VPWR),
    .Y(_03468_),
    .VSS(VGND),
    .A1(_03423_),
    .A2(_03421_));
 sg13g2_nand2_1 _09316_ (.Y(_03469_),
    .A(_03468_),
    .B(_03397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09317_ (.B1(_03469_),
    .VDD(VPWR),
    .Y(_03470_),
    .VSS(VGND),
    .A1(_03394_),
    .A2(_03392_));
 sg13g2_nand2_1 _09318_ (.Y(_03471_),
    .A(_03470_),
    .B(_03389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09319_ (.B1(_03471_),
    .VDD(VPWR),
    .Y(_03472_),
    .VSS(VGND),
    .A1(_03384_),
    .A2(_03386_));
 sg13g2_nand2_1 _09320_ (.Y(_03473_),
    .A(_03472_),
    .B(_03383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09321_ (.B1(_03473_),
    .VDD(VPWR),
    .Y(_03474_),
    .VSS(VGND),
    .A1(_03378_),
    .A2(_03380_));
 sg13g2_nand2_1 _09322_ (.Y(_03475_),
    .A(_03474_),
    .B(_03437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09323_ (.B1(_03475_),
    .VDD(VPWR),
    .Y(_03476_),
    .VSS(VGND),
    .A1(_03370_),
    .A2(_03434_));
 sg13g2_nand2_1 _09324_ (.Y(_03477_),
    .A(_03476_),
    .B(_03376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09325_ (.Y(_03478_),
    .A(\fp16_res_pipe.op_sign_logic0.mantisa_a[9] ),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _09326_ (.A2(_03478_),
    .A1(_03477_),
    .B1(_03446_),
    .X(_03479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09327_ (.B1(_03479_),
    .VDD(VPWR),
    .Y(_03480_),
    .VSS(VGND),
    .A1(_03444_),
    .A2(_03368_));
 sg13g2_nand2_1 _09328_ (.Y(_03481_),
    .A(_03480_),
    .B(_03365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09329_ (.Y(_03482_),
    .A(_03361_),
    .B(net1823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09330_ (.Y(_01276_),
    .A(_03481_),
    .B(_03482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09331_ (.B(_03446_),
    .C(_03478_),
    .A(_03477_),
    .Y(_03483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09332_ (.B(_03483_),
    .C(net1738),
    .A(_03479_),
    .Y(_03484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09333_ (.Y(_03485_),
    .A(net1770),
    .B(\fp16_res_pipe.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09334_ (.B1(_03375_),
    .VDD(VPWR),
    .Y(_03486_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.op_sign_logic0.mantisa_a[8] ),
    .A2(_03434_));
 sg13g2_inv_1 _09335_ (.VDD(VPWR),
    .Y(_03487_),
    .A(_03413_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09336_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03449_),
    .A2(_03415_),
    .Y(_03488_),
    .B1(_03487_));
 sg13g2_inv_1 _09337_ (.VDD(VPWR),
    .Y(_03489_),
    .A(_03488_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09338_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03489_),
    .A2(_03407_),
    .Y(_03490_),
    .B1(_03404_));
 sg13g2_a21oi_1 _09339_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03490_),
    .A2(_03418_),
    .Y(_03491_),
    .B1(_03401_));
 sg13g2_a21oi_1 _09340_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03491_),
    .A2(_03425_),
    .Y(_03492_),
    .B1(_03422_));
 sg13g2_a21oi_1 _09341_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03492_),
    .A2(_03428_),
    .Y(_03493_),
    .B1(_03395_));
 sg13g2_inv_1 _09342_ (.VDD(VPWR),
    .Y(_03494_),
    .A(_03493_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09343_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03382_),
    .A2(_03387_),
    .Y(_03495_),
    .B1(_03381_));
 sg13g2_o21ai_1 _09344_ (.B1(_03495_),
    .VDD(VPWR),
    .Y(_03496_),
    .VSS(VGND),
    .A1(_03391_),
    .A2(_03494_));
 sg13g2_a22oi_1 _09345_ (.Y(_03497_),
    .B1(_03438_),
    .B2(_03496_),
    .A2(_03486_),
    .A1(_03374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09346_ (.Y(_03498_),
    .A(_03440_),
    .B(_03452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09347_ (.B1(_03498_),
    .VDD(VPWR),
    .Y(_03499_),
    .VSS(VGND),
    .A1(_03445_),
    .A2(_03497_));
 sg13g2_inv_1 _09348_ (.VDD(VPWR),
    .Y(_03500_),
    .A(_03364_),
    .VSS(VGND));
 sg13g2_nor2_2 _09349_ (.A(_03361_),
    .B(_03500_),
    .Y(_03501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09350_ (.B(_03501_),
    .C(_03447_),
    .A(_03499_),
    .Y(_03502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09351_ (.B(_03485_),
    .C(_03502_),
    .A(_03484_),
    .Y(_01275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09352_ (.Y(_03503_),
    .B(_03377_),
    .A_N(_03476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09353_ (.B(net1738),
    .C(_03477_),
    .A(_03503_),
    .Y(_03504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09354_ (.Y(_03505_),
    .A(net1770),
    .B(\fp16_res_pipe.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09355_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03433_),
    .A2(_03436_),
    .Y(_03506_),
    .B1(_03371_));
 sg13g2_a21oi_1 _09356_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03496_),
    .A2(_03436_),
    .Y(_03507_),
    .B1(_03435_));
 sg13g2_nand2b_1 _09357_ (.Y(_03508_),
    .B(net1674),
    .A_N(_03507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09358_ (.B1(_03508_),
    .VDD(VPWR),
    .Y(_03509_),
    .VSS(VGND),
    .A1(net1674),
    .A2(_03506_));
 sg13g2_xnor2_1 _09359_ (.Y(_03510_),
    .A(_03376_),
    .B(_03509_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09360_ (.Y(_03511_),
    .A(_03510_),
    .B(_03501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09361_ (.B(_03505_),
    .C(_03511_),
    .A(_03504_),
    .Y(_01274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09362_ (.VDD(VPWR),
    .Y(_03512_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[8] ),
    .VSS(VGND));
 sg13g2_nand2b_1 _09363_ (.Y(_03513_),
    .B(net1674),
    .A_N(_03496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09364_ (.B1(_03513_),
    .VDD(VPWR),
    .Y(_03514_),
    .VSS(VGND),
    .A1(_03433_),
    .A2(net1674));
 sg13g2_xnor2_1 _09365_ (.Y(_03515_),
    .A(_03436_),
    .B(_03514_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09366_ (.A(_03437_),
    .B(_03474_),
    .Y(_03516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09367_ (.Y(_03517_),
    .A(_03475_),
    .B(\fp16_res_pipe.reg2en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _09368_ (.A(_03501_),
    .Y(_03518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09369_ (.B1(_03518_),
    .VDD(VPWR),
    .Y(_03519_),
    .VSS(VGND),
    .A1(_03516_),
    .A2(_03517_));
 sg13g2_o21ai_1 _09370_ (.B1(_03519_),
    .VDD(VPWR),
    .Y(_03520_),
    .VSS(VGND),
    .A1(_03500_),
    .A2(_03515_));
 sg13g2_o21ai_1 _09371_ (.B1(_03520_),
    .VDD(VPWR),
    .Y(_01273_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.reg2en.q[0] ),
    .A2(_03512_));
 sg13g2_a21oi_1 _09372_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03430_),
    .A2(_03388_),
    .Y(_03521_),
    .B1(_03385_));
 sg13g2_nor2_1 _09373_ (.A(_03389_),
    .B(_03494_),
    .Y(_03522_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09374_ (.B1(net1674),
    .VDD(VPWR),
    .Y(_03523_),
    .VSS(VGND),
    .A1(_03387_),
    .A2(_03522_));
 sg13g2_o21ai_1 _09375_ (.B1(_03523_),
    .VDD(VPWR),
    .Y(_03524_),
    .VSS(VGND),
    .A1(net1674),
    .A2(_03521_));
 sg13g2_xnor2_1 _09376_ (.Y(_03525_),
    .A(_03382_),
    .B(_03524_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09377_ (.Y(_03526_),
    .A(_03382_),
    .B(_03472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09378_ (.Y(_03527_),
    .B1(net1738),
    .B2(_03526_),
    .A2(\fp16_res_pipe.add_renorm0.mantisa[7] ),
    .A1(net1770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09379_ (.B1(_03527_),
    .VDD(VPWR),
    .Y(_01272_),
    .VSS(VGND),
    .A1(_03518_),
    .A2(_03525_));
 sg13g2_nand2_1 _09380_ (.Y(_03528_),
    .A(net1674),
    .B(_03493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09381_ (.B1(_03528_),
    .VDD(VPWR),
    .Y(_03529_),
    .VSS(VGND),
    .A1(_03431_),
    .A2(net1674));
 sg13g2_a21oi_1 _09382_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03529_),
    .A2(_03388_),
    .Y(_03530_),
    .B1(_03518_));
 sg13g2_o21ai_1 _09383_ (.B1(_03530_),
    .VDD(VPWR),
    .Y(_03531_),
    .VSS(VGND),
    .A1(_03388_),
    .A2(_03529_));
 sg13g2_nand2_1 _09384_ (.Y(_03532_),
    .A(net1770),
    .B(\fp16_res_pipe.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09385_ (.Y(_03533_),
    .B(_03388_),
    .A_N(_03470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09386_ (.B(net1738),
    .C(_03471_),
    .A(_03533_),
    .Y(_03534_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09387_ (.B(_03532_),
    .C(_03534_),
    .A(_03531_),
    .Y(_01271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03420_),
    .A2(_03425_),
    .Y(_03535_),
    .B1(_03424_));
 sg13g2_mux2_1 _09389_ (.A0(_03535_),
    .A1(_03492_),
    .S(net1675),
    .X(_03536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09390_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03536_),
    .A2(_03397_),
    .Y(_03537_),
    .B1(_03518_));
 sg13g2_o21ai_1 _09391_ (.B1(_03537_),
    .VDD(VPWR),
    .Y(_03538_),
    .VSS(VGND),
    .A1(_03397_),
    .A2(_03536_));
 sg13g2_inv_1 _09392_ (.VDD(VPWR),
    .Y(_03539_),
    .A(_03468_),
    .VSS(VGND));
 sg13g2_nand2_1 _09393_ (.Y(_03540_),
    .A(_03469_),
    .B(net1738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03396_),
    .A2(_03539_),
    .Y(_03541_),
    .B1(_03540_));
 sg13g2_a21oi_1 _09395_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1770),
    .A2(\fp16_res_pipe.add_renorm0.mantisa[5] ),
    .Y(_03542_),
    .B1(_03541_));
 sg13g2_nand2_1 _09396_ (.Y(_01270_),
    .A(_03538_),
    .B(_03542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _09397_ (.A0(_03420_),
    .A1(_03491_),
    .S(net1675),
    .X(_03543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09398_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03543_),
    .A2(_03425_),
    .Y(_03544_),
    .B1(_03518_));
 sg13g2_o21ai_1 _09399_ (.B1(_03544_),
    .VDD(VPWR),
    .Y(_03545_),
    .VSS(VGND),
    .A1(_03425_),
    .A2(_03543_));
 sg13g2_nand2_1 _09400_ (.Y(_03546_),
    .A(net1770),
    .B(\fp16_res_pipe.add_renorm0.mantisa[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09401_ (.Y(_03547_),
    .B(_03425_),
    .A_N(_03466_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09402_ (.B(net1738),
    .C(_03467_),
    .A(_03547_),
    .Y(_03548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09403_ (.B(_03546_),
    .C(_03548_),
    .A(_03545_),
    .Y(_01269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09404_ (.VDD(VPWR),
    .Y(_03549_),
    .A(_03406_),
    .VSS(VGND));
 sg13g2_o21ai_1 _09405_ (.B1(_03549_),
    .VDD(VPWR),
    .Y(_03550_),
    .VSS(VGND),
    .A1(_03404_),
    .A2(_03417_));
 sg13g2_nand2_1 _09406_ (.Y(_03551_),
    .A(net1675),
    .B(_03490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09407_ (.B1(_03551_),
    .VDD(VPWR),
    .Y(_03552_),
    .VSS(VGND),
    .A1(net1675),
    .A2(_03550_));
 sg13g2_a21oi_1 _09408_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03552_),
    .A2(_03464_),
    .Y(_03553_),
    .B1(_03518_));
 sg13g2_o21ai_1 _09409_ (.B1(_03553_),
    .VDD(VPWR),
    .Y(_03554_),
    .VSS(VGND),
    .A1(_03464_),
    .A2(_03552_));
 sg13g2_nand2_1 _09410_ (.Y(_03555_),
    .A(_03361_),
    .B(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09411_ (.Y(_03556_),
    .B(_03402_),
    .A_N(_03463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09412_ (.B(net1738),
    .C(_03465_),
    .A(_03556_),
    .Y(_03557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09413_ (.B(_03555_),
    .C(_03557_),
    .A(_03554_),
    .Y(_01268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09414_ (.Y(_03558_),
    .A(net1675),
    .B(_03489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09415_ (.B1(_03558_),
    .VDD(VPWR),
    .Y(_03559_),
    .VSS(VGND),
    .A1(_03417_),
    .A2(net1675));
 sg13g2_and2_1 _09416_ (.A(_03559_),
    .B(_03407_),
    .X(_03560_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09417_ (.B1(_03501_),
    .VDD(VPWR),
    .Y(_03561_),
    .VSS(VGND),
    .A1(_03407_),
    .A2(_03559_));
 sg13g2_nand2b_1 _09418_ (.Y(_03562_),
    .B(_03407_),
    .A_N(_03461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _09419_ (.A(_03462_),
    .B(net1738),
    .X(_03563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09420_ (.Y(_03564_),
    .B1(_03562_),
    .B2(_03563_),
    .A2(\fp16_res_pipe.add_renorm0.mantisa[2] ),
    .A1(net1770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09421_ (.B1(_03564_),
    .VDD(VPWR),
    .Y(_01267_),
    .VSS(VGND),
    .A1(_03560_),
    .A2(_03561_));
 sg13g2_inv_1 _09422_ (.VDD(VPWR),
    .Y(_03565_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[1] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _09423_ (.Y(_03566_),
    .A(_03459_),
    .B(_03443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09424_ (.Y(_03567_),
    .A(net1675),
    .B(_03449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09425_ (.B1(_03567_),
    .VDD(VPWR),
    .Y(_03568_),
    .VSS(VGND),
    .A1(_03410_),
    .A2(net1675));
 sg13g2_xor2_1 _09426_ (.B(_03568_),
    .A(_03443_),
    .X(_03569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09427_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03569_),
    .A2(_03364_),
    .Y(_03570_),
    .B1(net1770));
 sg13g2_o21ai_1 _09428_ (.B1(_03570_),
    .VDD(VPWR),
    .Y(_03571_),
    .VSS(VGND),
    .A1(_03364_),
    .A2(_03566_));
 sg13g2_o21ai_1 _09429_ (.B1(_03571_),
    .VDD(VPWR),
    .Y(_01266_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.reg2en.q[0] ),
    .A2(_03565_));
 sg13g2_inv_1 _09430_ (.VDD(VPWR),
    .Y(_03572_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09431_ (.Y(_03573_),
    .A(_03450_),
    .B(\fp16_res_pipe.reg2en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09432_ (.B1(_03573_),
    .VDD(VPWR),
    .Y(_01265_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.reg2en.q[0] ),
    .A2(_03572_));
 sg13g2_inv_1 _09433_ (.VDD(VPWR),
    .Y(_03574_),
    .A(\fp16_res_pipe.add_renorm0.exp[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09434_ (.Y(_03575_),
    .A(net1833),
    .B(\fp16_res_pipe.seg_reg0.q[29] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09435_ (.B1(_03575_),
    .VDD(VPWR),
    .Y(_01264_),
    .VSS(VGND),
    .A1(net1834),
    .A2(_03574_));
 sg13g2_inv_2 _09436_ (.Y(_03576_),
    .A(\fp16_res_pipe.add_renorm0.exp[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09437_ (.Y(_03577_),
    .A(net1834),
    .B(\fp16_res_pipe.seg_reg0.q[28] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09438_ (.B1(_03577_),
    .VDD(VPWR),
    .Y(_01263_),
    .VSS(VGND),
    .A1(net1834),
    .A2(_03576_));
 sg13g2_inv_1 _09439_ (.VDD(VPWR),
    .Y(_03578_),
    .A(\fp16_res_pipe.add_renorm0.exp[5] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09440_ (.Y(_03579_),
    .A(net1834),
    .B(\fp16_res_pipe.seg_reg0.q[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09441_ (.B1(_03579_),
    .VDD(VPWR),
    .Y(_01262_),
    .VSS(VGND),
    .A1(net1834),
    .A2(_03578_));
 sg13g2_inv_2 _09442_ (.Y(_03580_),
    .A(\fp16_res_pipe.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09443_ (.Y(_03581_),
    .A(net1833),
    .B(\fp16_res_pipe.seg_reg0.q[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09444_ (.B1(_03581_),
    .VDD(VPWR),
    .Y(_01261_),
    .VSS(VGND),
    .A1(net1832),
    .A2(_03580_));
 sg13g2_inv_1 _09445_ (.VDD(VPWR),
    .Y(_03582_),
    .A(\fp16_res_pipe.add_renorm0.exp[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09446_ (.Y(_03583_),
    .A(net1833),
    .B(\fp16_res_pipe.seg_reg0.q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09447_ (.B1(_03583_),
    .VDD(VPWR),
    .Y(_01260_),
    .VSS(VGND),
    .A1(net1832),
    .A2(_03582_));
 sg13g2_inv_1 _09448_ (.VDD(VPWR),
    .Y(_03584_),
    .A(\fp16_res_pipe.add_renorm0.exp[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09449_ (.Y(_03585_),
    .A(net1832),
    .B(\fp16_res_pipe.seg_reg0.q[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09450_ (.B1(_03585_),
    .VDD(VPWR),
    .Y(_01259_),
    .VSS(VGND),
    .A1(net1832),
    .A2(_03584_));
 sg13g2_inv_2 _09451_ (.Y(_03586_),
    .A(\fp16_res_pipe.add_renorm0.exp[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09452_ (.Y(_03587_),
    .A(net1832),
    .B(\fp16_res_pipe.seg_reg0.q[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09453_ (.B1(_03587_),
    .VDD(VPWR),
    .Y(_01258_),
    .VSS(VGND),
    .A1(net1832),
    .A2(_03586_));
 sg13g2_mux2_1 _09454_ (.A0(\fp16_res_pipe.add_renorm0.exp[0] ),
    .A1(\fp16_res_pipe.seg_reg0.q[22] ),
    .S(net1833),
    .X(_01257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09455_ (.A(\fp16_res_pipe.exp_mant_logic0.a[15] ),
    .B(net1911),
    .Y(_03588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09456_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03327_),
    .A2(net1911),
    .Y(_01256_),
    .B1(_03588_));
 sg13g2_inv_1 _09457_ (.VDD(VPWR),
    .Y(_03589_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[14] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09458_ (.Y(_03590_),
    .A(\acc_sub.x2[14] ),
    .B(net1915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09459_ (.B1(_03590_),
    .VDD(VPWR),
    .Y(_01255_),
    .VSS(VGND),
    .A1(net1915),
    .A2(_03589_));
 sg13g2_inv_1 _09460_ (.VDD(VPWR),
    .Y(_03591_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[13] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09461_ (.Y(_03592_),
    .A(\acc_sub.x2[13] ),
    .B(net1915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09462_ (.B1(_03592_),
    .VDD(VPWR),
    .Y(_01254_),
    .VSS(VGND),
    .A1(net1915),
    .A2(_03591_));
 sg13g2_inv_1 _09463_ (.VDD(VPWR),
    .Y(_03593_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09464_ (.Y(_03594_),
    .A(\acc_sub.x2[12] ),
    .B(net1913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09465_ (.B1(_03594_),
    .VDD(VPWR),
    .Y(_01253_),
    .VSS(VGND),
    .A1(net1915),
    .A2(_03593_));
 sg13g2_inv_1 _09466_ (.VDD(VPWR),
    .Y(_03595_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09467_ (.Y(_03596_),
    .A(\acc_sub.x2[11] ),
    .B(net1914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09468_ (.B1(_03596_),
    .VDD(VPWR),
    .Y(_01252_),
    .VSS(VGND),
    .A1(net1914),
    .A2(_03595_));
 sg13g2_inv_1 _09469_ (.VDD(VPWR),
    .Y(_03597_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09470_ (.Y(_03598_),
    .A(\acc_sub.x2[10] ),
    .B(net1914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09471_ (.B1(_03598_),
    .VDD(VPWR),
    .Y(_01251_),
    .VSS(VGND),
    .A1(net1914),
    .A2(_03597_));
 sg13g2_inv_1 _09472_ (.VDD(VPWR),
    .Y(_03599_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09473_ (.Y(_03600_),
    .A(\acc_sub.x2[9] ),
    .B(net1912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09474_ (.B1(_03600_),
    .VDD(VPWR),
    .Y(_01250_),
    .VSS(VGND),
    .A1(net1920),
    .A2(_03599_));
 sg13g2_inv_4 _09475_ (.A(\acc_sub.x2[8] ),
    .Y(_03601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09476_ (.A(net1919),
    .B(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .Y(_03602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09477_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03601_),
    .A2(net1919),
    .Y(_01249_),
    .B1(_03602_));
 sg13g2_inv_4 _09478_ (.A(\acc_sub.x2[7] ),
    .Y(_03603_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09479_ (.A(net1919),
    .B(\fp16_res_pipe.exp_mant_logic0.a[7] ),
    .Y(_03604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03603_),
    .A2(net1919),
    .Y(_01248_),
    .B1(_03604_));
 sg13g2_inv_2 _09481_ (.Y(_03605_),
    .A(net1827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09482_ (.Y(_03606_),
    .A(\acc_sub.x2[6] ),
    .B(net1916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09483_ (.B1(_03606_),
    .VDD(VPWR),
    .Y(_01247_),
    .VSS(VGND),
    .A1(net1917),
    .A2(_03605_));
 sg13g2_inv_2 _09484_ (.Y(_03607_),
    .A(net1828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09485_ (.Y(_03608_),
    .A(\acc_sub.x2[5] ),
    .B(net1917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09486_ (.B1(_03608_),
    .VDD(VPWR),
    .Y(_01246_),
    .VSS(VGND),
    .A1(net1917),
    .A2(_03607_));
 sg13g2_inv_2 _09487_ (.Y(_03609_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09488_ (.Y(_03610_),
    .A(\acc_sub.x2[4] ),
    .B(net1918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09489_ (.B1(_03610_),
    .VDD(VPWR),
    .Y(_01245_),
    .VSS(VGND),
    .A1(net1918),
    .A2(_03609_));
 sg13g2_inv_2 _09490_ (.Y(_03611_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09491_ (.Y(_03612_),
    .A(\acc_sub.x2[3] ),
    .B(net1918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09492_ (.B1(_03612_),
    .VDD(VPWR),
    .Y(_01244_),
    .VSS(VGND),
    .A1(net1918),
    .A2(_03611_));
 sg13g2_inv_2 _09493_ (.Y(_03613_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09494_ (.Y(_03614_),
    .A(\acc_sub.x2[2] ),
    .B(net1918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09495_ (.B1(_03614_),
    .VDD(VPWR),
    .Y(_01243_),
    .VSS(VGND),
    .A1(net1917),
    .A2(_03613_));
 sg13g2_inv_2 _09496_ (.Y(_03615_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09497_ (.Y(_03616_),
    .A(\acc_sub.x2[1] ),
    .B(net1916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09498_ (.B1(_03616_),
    .VDD(VPWR),
    .Y(_01242_),
    .VSS(VGND),
    .A1(net1916),
    .A2(_03615_));
 sg13g2_inv_2 _09499_ (.Y(_03617_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09500_ (.Y(_03618_),
    .A(\acc_sub.x2[0] ),
    .B(net1916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09501_ (.B1(_03618_),
    .VDD(VPWR),
    .Y(_01241_),
    .VSS(VGND),
    .A1(net1916),
    .A2(_03617_));
 sg13g2_inv_1 _09502_ (.VDD(VPWR),
    .Y(_03619_),
    .A(\acc_sum.add_renorm0.mantisa[9] ),
    .VSS(VGND));
 sg13g2_inv_1 _09503_ (.VDD(VPWR),
    .Y(_03620_),
    .A(\acc_sum.add_renorm0.mantisa[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09504_ (.Y(_03621_),
    .A(\acc_sum.add_renorm0.mantisa[3] ),
    .B(\acc_sum.add_renorm0.mantisa[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09505_ (.VDD(VPWR),
    .Y(_03622_),
    .A(_03621_),
    .VSS(VGND));
 sg13g2_nand3_1 _09506_ (.B(\acc_sum.add_renorm0.mantisa[5] ),
    .C(\acc_sum.add_renorm0.mantisa[4] ),
    .A(_03622_),
    .Y(_03623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09507_ (.A(_03620_),
    .B(_03623_),
    .Y(_03624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09508_ (.B(\acc_sum.add_renorm0.mantisa[8] ),
    .C(\acc_sum.add_renorm0.mantisa[7] ),
    .A(_03624_),
    .Y(_03625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1755 (.A(_06750_),
    .X(net1755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09510_ (.A(_03619_),
    .B(_03625_),
    .Y(_03627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09511_ (.A(\acc_sum.add_renorm0.mantisa[10] ),
    .B(_03627_),
    .Y(_03628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1707 (.A(_02652_),
    .X(net1707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _09513_ (.A(_03628_),
    .Y(_03630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09514_ (.Y(_03631_),
    .A(\acc_sum.add_renorm0.mantisa[6] ),
    .B(_03623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout94 (.A(net96),
    .X(net94),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09516_ (.Y(_03633_),
    .A(_03631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09517_ (.Y(_03634_),
    .A(\acc_sum.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09518_ (.Y(_03635_),
    .A(_03634_),
    .B(_03624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1759 (.A(_04993_),
    .X(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09520_ (.VDD(VPWR),
    .Y(_03637_),
    .A(_03624_),
    .VSS(VGND));
 sg13g2_inv_1 _09521_ (.VDD(VPWR),
    .Y(_03638_),
    .A(\acc_sum.add_renorm0.mantisa[8] ),
    .VSS(VGND));
 sg13g2_o21ai_1 _09522_ (.B1(_03638_),
    .VDD(VPWR),
    .Y(_03639_),
    .VSS(VGND),
    .A1(_03634_),
    .A2(_03637_));
 sg13g2_nand2_2 _09523_ (.Y(_03640_),
    .A(_03639_),
    .B(_03625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09524_ (.VDD(VPWR),
    .Y(_03641_),
    .A(_03640_),
    .VSS(VGND));
 sg13g2_inv_1 _09525_ (.VDD(VPWR),
    .Y(_03642_),
    .A(_03627_),
    .VSS(VGND));
 sg13g2_nand2_1 _09526_ (.Y(_03643_),
    .A(_03625_),
    .B(_03619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09527_ (.Y(_03644_),
    .A(_03642_),
    .B(_03643_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09528_ (.VDD(VPWR),
    .Y(_03645_),
    .A(_03644_),
    .VSS(VGND));
 sg13g2_nor4_1 _09529_ (.A(_03633_),
    .B(_03635_),
    .C(_03641_),
    .D(_03645_),
    .Y(_03646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09530_ (.A(_03630_),
    .B(_03646_),
    .Y(_03647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09531_ (.Y(_03648_),
    .A(_03647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _09532_ (.A(_03640_),
    .B(_03630_),
    .C(_03645_),
    .Y(_03649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09533_ (.VDD(VPWR),
    .Y(_03650_),
    .A(\acc_sum.add_renorm0.mantisa[5] ),
    .VSS(VGND));
 sg13g2_nor2b_1 _09534_ (.A(_03621_),
    .B_N(\acc_sum.add_renorm0.mantisa[4] ),
    .Y(_03651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09535_ (.Y(_03652_),
    .A(_03650_),
    .B(_03651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout82 (.A(net83),
    .X(net82),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09537_ (.VDD(VPWR),
    .Y(_03654_),
    .A(_03652_),
    .VSS(VGND));
 sg13g2_xnor2_1 _09538_ (.Y(_03655_),
    .A(\acc_sum.add_renorm0.mantisa[4] ),
    .B(_03621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout65 (.A(net66),
    .X(net65),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09540_ (.B(_03654_),
    .C(_03655_),
    .A(_03633_),
    .Y(_03657_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09541_ (.B(_03628_),
    .C(_03640_),
    .A(_03644_),
    .Y(_03658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09542_ (.A(_03635_),
    .B(_03658_),
    .Y(_03659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09543_ (.VDD(VPWR),
    .Y(_03660_),
    .A(_03659_),
    .VSS(VGND));
 sg13g2_nor2_2 _09544_ (.A(_03657_),
    .B(_03660_),
    .Y(_03661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09545_ (.A(_03649_),
    .B(_03661_),
    .Y(_03662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _09546_ (.A(_03662_),
    .Y(_03663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09547_ (.A(_03648_),
    .B(_03663_),
    .Y(_03664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09548_ (.VDD(VPWR),
    .Y(_03665_),
    .A(_03664_),
    .VSS(VGND));
 sg13g2_nor2_2 _09549_ (.A(_03644_),
    .B(_03630_),
    .Y(_03666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _09550_ (.X(_03667_),
    .A(_03659_),
    .B(_03652_),
    .C(_03633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1689 (.A(_04050_),
    .X(net1689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09552_ (.VDD(VPWR),
    .Y(_03669_),
    .A(\acc_sum.add_renorm0.mantisa[1] ),
    .VSS(VGND));
 sg13g2_inv_1 _09553_ (.VDD(VPWR),
    .Y(_03670_),
    .A(\acc_sum.add_renorm0.mantisa[2] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _09554_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03669_),
    .A2(_02918_),
    .Y(_03671_),
    .B1(_03670_));
 sg13g2_inv_1 _09555_ (.VDD(VPWR),
    .Y(_03672_),
    .A(_03671_),
    .VSS(VGND));
 sg13g2_inv_2 _09556_ (.Y(_03673_),
    .A(\acc_sum.add_renorm0.mantisa[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09557_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03622_),
    .Y(_03674_),
    .A2(_03673_),
    .A1(_03672_));
 sg13g2_inv_1 _09558_ (.VDD(VPWR),
    .Y(_03675_),
    .A(_03674_),
    .VSS(VGND));
 sg13g2_nor4_1 _09559_ (.A(_03652_),
    .B(_03655_),
    .C(_03675_),
    .D(_03631_),
    .Y(_03676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09560_ (.Y(_03677_),
    .A(_03659_),
    .B(_03676_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _09561_ (.A(_03667_),
    .B_N(_03677_),
    .Y(_03678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09562_ (.VDD(VPWR),
    .Y(_03679_),
    .A(_03658_),
    .VSS(VGND));
 sg13g2_nand2_2 _09563_ (.Y(_03680_),
    .A(_03679_),
    .B(_03635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _09564_ (.B(_03678_),
    .C(_03680_),
    .Y(_03681_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_03666_));
 sg13g2_buf_2 place1671 (.A(_02800_),
    .X(net1671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09566_ (.B1(net1803),
    .VDD(VPWR),
    .Y(_03683_),
    .VSS(VGND),
    .A1(_03665_),
    .A2(_03681_));
 sg13g2_nor2_2 _09567_ (.A(_03633_),
    .B(_03660_),
    .Y(_03684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09568_ (.Y(_03685_),
    .B1(_03674_),
    .B2(_03667_),
    .A2(_03684_),
    .A1(_03655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09569_ (.Y(_03686_),
    .B1(_03635_),
    .B2(_03666_),
    .A2(_03641_),
    .A1(_03630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09570_ (.VDD(VPWR),
    .Y(_03687_),
    .A(_03680_),
    .VSS(VGND));
 sg13g2_a22oi_1 _09571_ (.Y(_03688_),
    .B1(_03652_),
    .B2(_03687_),
    .A2(_03649_),
    .A1(_03631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09572_ (.B(_03686_),
    .C(_03688_),
    .A(_03685_),
    .Y(_03689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09573_ (.Y(_03690_),
    .A(net1806),
    .B(\acc_sum.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09574_ (.B1(_03690_),
    .VDD(VPWR),
    .Y(_03691_),
    .VSS(VGND),
    .A1(net1806),
    .A2(_03620_));
 sg13g2_inv_1 _09575_ (.VDD(VPWR),
    .Y(_03692_),
    .A(_03691_),
    .VSS(VGND));
 sg13g2_nand2_1 _09576_ (.Y(_03693_),
    .A(net1806),
    .B(\acc_sum.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09577_ (.B1(_03693_),
    .VDD(VPWR),
    .Y(_03694_),
    .VSS(VGND),
    .A1(net1806),
    .A2(_03638_));
 sg13g2_nand2_1 _09578_ (.Y(_03695_),
    .A(net1806),
    .B(\acc_sum.add_renorm0.mantisa[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09579_ (.B1(_03695_),
    .VDD(VPWR),
    .Y(_03696_),
    .VSS(VGND),
    .A1(net1806),
    .A2(_03634_));
 sg13g2_nand2_1 _09580_ (.Y(_03697_),
    .A(_03694_),
    .B(_03696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09581_ (.Y(_03698_),
    .A(net1805),
    .B(\acc_sum.add_renorm0.mantisa[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09582_ (.VDD(VPWR),
    .Y(_03699_),
    .A(_03698_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09583_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_02806_),
    .A2(\acc_sum.add_renorm0.mantisa[4] ),
    .Y(_03700_),
    .B1(_03699_));
 sg13g2_inv_1 _09584_ (.VDD(VPWR),
    .Y(_03701_),
    .A(_03700_),
    .VSS(VGND));
 sg13g2_nand2_1 _09585_ (.Y(_03702_),
    .A(_02806_),
    .B(_03673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09586_ (.B1(_03702_),
    .VDD(VPWR),
    .Y(_03703_),
    .VSS(VGND),
    .A1(_02806_),
    .A2(\acc_sum.add_renorm0.mantisa[4] ));
 sg13g2_inv_1 _09587_ (.VDD(VPWR),
    .Y(_03704_),
    .A(_03703_),
    .VSS(VGND));
 sg13g2_nand2_1 _09588_ (.Y(_03705_),
    .A(net1805),
    .B(\acc_sum.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09589_ (.B1(_03705_),
    .VDD(VPWR),
    .Y(_03706_),
    .VSS(VGND),
    .A1(net1805),
    .A2(_03650_));
 sg13g2_nand3_1 _09590_ (.B(_03704_),
    .C(_03706_),
    .A(_03701_),
    .Y(_03707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09591_ (.A(net1805),
    .B(\acc_sum.add_renorm0.mantisa[2] ),
    .Y(_03708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09592_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1805),
    .A2(_03673_),
    .Y(_03709_),
    .B1(_03708_));
 sg13g2_inv_2 _09593_ (.Y(_03710_),
    .A(_03709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09594_ (.A(_03703_),
    .B(_03710_),
    .Y(_03711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09595_ (.Y(_03712_),
    .B1(_02806_),
    .B2(_02918_),
    .A2(\acc_sum.add_renorm0.mantisa[3] ),
    .A1(_03670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _09596_ (.A(\acc_sum.add_renorm0.mantisa[1] ),
    .B(_03708_),
    .C(_03712_),
    .Y(_03713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09597_ (.A(_03710_),
    .B(_03713_),
    .Y(_03714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09598_ (.A(_03711_),
    .B(_03714_),
    .Y(_03715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09599_ (.A(_03707_),
    .B(_03715_),
    .Y(_03716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09600_ (.VDD(VPWR),
    .Y(_03717_),
    .A(_03716_),
    .VSS(VGND));
 sg13g2_nor3_1 _09601_ (.A(_03692_),
    .B(_03697_),
    .C(_03717_),
    .Y(_03718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09602_ (.A(_03692_),
    .B(_03717_),
    .Y(_03719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03719_),
    .A2(_03696_),
    .Y(_03720_),
    .B1(_03694_));
 sg13g2_nor3_1 _09604_ (.A(net1804),
    .B(_03718_),
    .C(_03720_),
    .Y(_03721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09605_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03689_),
    .A2(net1804),
    .Y(_03722_),
    .B1(_03721_));
 sg13g2_nor2_2 _09606_ (.A(net1805),
    .B(\acc_sum.add_renorm0.mantisa[10] ),
    .Y(_03723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09607_ (.Y(_03724_),
    .A(net1806),
    .B(\acc_sum.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09608_ (.B1(_03724_),
    .VDD(VPWR),
    .Y(_03725_),
    .VSS(VGND),
    .A1(net1805),
    .A2(_03619_));
 sg13g2_inv_1 _09609_ (.VDD(VPWR),
    .Y(_03726_),
    .A(_03725_),
    .VSS(VGND));
 sg13g2_nor2_1 _09610_ (.A(_03692_),
    .B(_03697_),
    .Y(_03727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09611_ (.Y(_03728_),
    .B(_03727_),
    .A_N(_03707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09612_ (.A(_03726_),
    .B(_03728_),
    .Y(_03729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09613_ (.VDD(VPWR),
    .Y(_03730_),
    .A(_03729_),
    .VSS(VGND));
 sg13g2_nor2_1 _09614_ (.A(_03723_),
    .B(_03730_),
    .Y(_03731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09615_ (.VDD(VPWR),
    .Y(_03732_),
    .A(_03715_),
    .VSS(VGND));
 sg13g2_nand2_1 _09616_ (.Y(_03733_),
    .A(_03731_),
    .B(_03732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09617_ (.VDD(VPWR),
    .Y(_03734_),
    .A(_03733_),
    .VSS(VGND));
 sg13g2_xnor2_1 _09618_ (.Y(_03735_),
    .A(_03723_),
    .B(_03729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09619_ (.Y(_03736_),
    .A(_03735_),
    .B(_03713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09620_ (.Y(_03737_),
    .A(_03735_),
    .B(_03714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09621_ (.Y(_03738_),
    .B(_03710_),
    .A_N(_03723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09622_ (.B(_03737_),
    .C(_03738_),
    .A(_03736_),
    .Y(_03739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _09623_ (.A(net1802),
    .Y(_03740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09624_ (.B1(_03740_),
    .VDD(VPWR),
    .Y(_03741_),
    .VSS(VGND),
    .A1(_03734_),
    .A2(_03739_));
 sg13g2_xnor2_1 _09625_ (.Y(_03742_),
    .A(_03696_),
    .B(_03719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09626_ (.A(net1802),
    .B(_03742_),
    .Y(_03743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09627_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03704_),
    .A2(_03710_),
    .Y(_03744_),
    .B1(_03714_));
 sg13g2_a21oi_1 _09628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03704_),
    .A2(_03714_),
    .Y(_03745_),
    .B1(_03744_));
 sg13g2_o21ai_1 _09629_ (.B1(net1804),
    .VDD(VPWR),
    .Y(_03746_),
    .VSS(VGND),
    .A1(_03675_),
    .A2(_03628_));
 sg13g2_o21ai_1 _09630_ (.B1(_03746_),
    .VDD(VPWR),
    .Y(_03747_),
    .VSS(VGND),
    .A1(\acc_sum.seg_reg1.q[21] ),
    .A2(_03745_));
 sg13g2_nor2b_1 _09631_ (.A(_03743_),
    .B_N(_03747_),
    .Y(_03748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _09632_ (.A(_03683_),
    .B(_03722_),
    .C(_03741_),
    .D(_03748_),
    .X(_03749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09633_ (.Y(_03750_),
    .A(_03691_),
    .B(_03716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09634_ (.A(_03675_),
    .B(_03680_),
    .Y(_03751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09635_ (.Y(_03752_),
    .A(_03649_),
    .B(_03655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09636_ (.Y(_03753_),
    .A(_03666_),
    .B(_03652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09637_ (.Y(_03754_),
    .A(_03630_),
    .B(_03631_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09638_ (.B(_03753_),
    .C(_03754_),
    .A(_03752_),
    .Y(_03755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09639_ (.B1(net1804),
    .VDD(VPWR),
    .Y(_03756_),
    .VSS(VGND),
    .A1(_03751_),
    .A2(_03755_));
 sg13g2_o21ai_1 _09640_ (.B1(_03756_),
    .VDD(VPWR),
    .Y(_03757_),
    .VSS(VGND),
    .A1(net1802),
    .A2(_03750_));
 sg13g2_a21oi_1 _09641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03711_),
    .A2(_03701_),
    .Y(_03758_),
    .B1(_03706_));
 sg13g2_nand2b_1 _09642_ (.Y(_03759_),
    .B(_03717_),
    .A_N(_03758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09643_ (.Y(_03760_),
    .A(_03649_),
    .B(_03674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09644_ (.Y(_03761_),
    .A(_03630_),
    .B(_03652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09645_ (.Y(_03762_),
    .A(_03666_),
    .B(_03655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09646_ (.B(_03761_),
    .C(_03762_),
    .A(_03760_),
    .Y(_03763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09647_ (.Y(_03764_),
    .A(_03763_),
    .B(net1802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09648_ (.B1(_03764_),
    .VDD(VPWR),
    .Y(_03765_),
    .VSS(VGND),
    .A1(net1802),
    .A2(_03759_));
 sg13g2_a22oi_1 _09649_ (.Y(_03766_),
    .B1(_03655_),
    .B2(_03667_),
    .A2(_03684_),
    .A1(_03652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09650_ (.Y(_03767_),
    .A(_03628_),
    .B(_03640_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09651_ (.Y(_03768_),
    .B1(_03631_),
    .B2(_03687_),
    .A2(_03767_),
    .A1(_03645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09652_ (.Y(_03769_),
    .B1(_03674_),
    .B2(_03661_),
    .A2(_03649_),
    .A1(_03635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09653_ (.B(_03768_),
    .C(_03769_),
    .A(_03766_),
    .Y(_03770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09654_ (.Y(_03771_),
    .A(_03728_),
    .B(_03726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09655_ (.B(_03732_),
    .C(_03771_),
    .A(_03730_),
    .Y(_03772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09656_ (.B1(_03772_),
    .VDD(VPWR),
    .Y(_03773_),
    .VSS(VGND),
    .A1(_03732_),
    .A2(_03726_));
 sg13g2_and2_1 _09657_ (.A(_03773_),
    .B(_03740_),
    .X(_03774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09658_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03774_),
    .Y(_03775_),
    .A2(net1802),
    .A1(_03770_));
 sg13g2_xnor2_1 _09659_ (.Y(_03776_),
    .A(_03700_),
    .B(_03711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09660_ (.Y(_03777_),
    .B1(_03674_),
    .B2(_03666_),
    .A2(_03655_),
    .A1(_03630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09661_ (.A(_03740_),
    .B(_03777_),
    .Y(_03778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09662_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03778_),
    .Y(_03779_),
    .A2(_03776_),
    .A1(_03740_));
 sg13g2_nand2_1 _09663_ (.Y(_03780_),
    .A(_03775_),
    .B(_03779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _09664_ (.A(_03757_),
    .B(_03765_),
    .C(_03780_),
    .Y(_03781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09665_ (.Y(_03782_),
    .A(\acc_sum.reg3en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09666_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03782_),
    .Y(_03783_),
    .A2(_03781_),
    .A1(_03749_));
 sg13g2_buf_2 place1649 (.A(_01959_),
    .X(net1649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09668_ (.VDD(VPWR),
    .Y(_03785_),
    .A(_03783_),
    .VSS(VGND));
 sg13g2_buf_2 fanout51 (.A(net56),
    .X(net51),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09670_ (.Y(_03787_),
    .A(_03782_),
    .B(\acc_sum.y[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09671_ (.B1(_03787_),
    .VDD(VPWR),
    .Y(_01240_),
    .VSS(VGND),
    .A1(_02729_),
    .A2(_03785_));
 sg13g2_nand3_1 _09672_ (.B(\acc_sum.add_renorm0.exp[1] ),
    .C(\acc_sum.add_renorm0.exp[0] ),
    .A(\acc_sum.add_renorm0.exp[2] ),
    .Y(_03788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09673_ (.A(_02926_),
    .B(_03788_),
    .Y(_03789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09674_ (.Y(_03790_),
    .A(_03789_),
    .B(\acc_sum.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09675_ (.A(_02924_),
    .B(_03790_),
    .Y(_03791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09676_ (.Y(_03792_),
    .A(_03791_),
    .B(\acc_sum.add_renorm0.exp[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09677_ (.Y(_03793_),
    .A(_02920_),
    .B(_03792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09678_ (.A(net1807),
    .B(\acc_sum.add_renorm0.exp[7] ),
    .Y(_03794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09679_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03793_),
    .A2(net1807),
    .Y(_03795_),
    .B1(_03794_));
 sg13g2_xnor2_1 _09680_ (.Y(_03796_),
    .A(\acc_sum.add_renorm0.exp[5] ),
    .B(_03790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09681_ (.Y(_03797_),
    .A(_03796_),
    .B(net1807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09682_ (.B1(_03797_),
    .VDD(VPWR),
    .Y(_03798_),
    .VSS(VGND),
    .A1(net1807),
    .A2(_02924_));
 sg13g2_inv_1 _09683_ (.VDD(VPWR),
    .Y(_03799_),
    .A(_03798_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09684_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc_sum.add_renorm0.exp[1] ),
    .A2(\acc_sum.add_renorm0.exp[0] ),
    .Y(_03800_),
    .B1(\acc_sum.add_renorm0.exp[2] ));
 sg13g2_nor2b_1 _09685_ (.A(_03800_),
    .B_N(_03788_),
    .Y(_03801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09686_ (.Y(_03802_),
    .A(_03801_),
    .B(\acc_sum.add_renorm0.mantisa[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09687_ (.B1(_03802_),
    .VDD(VPWR),
    .Y(_03803_),
    .VSS(VGND),
    .A1(\acc_sum.add_renorm0.mantisa[11] ),
    .A2(_02928_));
 sg13g2_inv_1 _09688_ (.VDD(VPWR),
    .Y(_03804_),
    .A(_03803_),
    .VSS(VGND));
 sg13g2_nor2_1 _09689_ (.A(\acc_sum.add_renorm0.mantisa[11] ),
    .B(\acc_sum.add_renorm0.exp[0] ),
    .Y(_03805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09690_ (.Y(_03806_),
    .A(\acc_sum.add_renorm0.mantisa[11] ),
    .B(\acc_sum.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _09691_ (.A(_03805_),
    .B_N(_03806_),
    .Y(_03807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09692_ (.B(\acc_sum.add_renorm0.exp[1] ),
    .C(_03807_),
    .A(_03734_),
    .Y(_03808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09693_ (.A(_03804_),
    .B(_03808_),
    .Y(_03809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09694_ (.Y(_03810_),
    .A(_02926_),
    .B(_03788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09695_ (.Y(_03811_),
    .A(_02806_),
    .B(\acc_sum.add_renorm0.exp[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09696_ (.B1(_03811_),
    .VDD(VPWR),
    .Y(_03812_),
    .VSS(VGND),
    .A1(_02806_),
    .A2(_03810_));
 sg13g2_and2_1 _09697_ (.A(_03809_),
    .B(_03812_),
    .X(_03813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1672 (.A(_01847_),
    .X(net1672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09699_ (.Y(_03815_),
    .A(\acc_sum.add_renorm0.exp[4] ),
    .B(_03789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09700_ (.A(net1807),
    .B(\acc_sum.add_renorm0.exp[4] ),
    .Y(_03816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09701_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03815_),
    .A2(net1807),
    .Y(_03817_),
    .B1(_03816_));
 sg13g2_nand2_1 _09702_ (.Y(_03818_),
    .A(_03813_),
    .B(_03817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09703_ (.A(_03799_),
    .B(_03818_),
    .Y(_03819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09704_ (.Y(_03820_),
    .A(\acc_sum.add_renorm0.exp[6] ),
    .B(_03791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09705_ (.A(net1807),
    .B(\acc_sum.add_renorm0.exp[6] ),
    .Y(_03821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09706_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03820_),
    .A2(net1807),
    .Y(_03822_),
    .B1(_03821_));
 sg13g2_nand2_1 _09707_ (.Y(_03823_),
    .A(_03819_),
    .B(_03822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1790 (.A(net1788),
    .X(net1790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09709_ (.B1(net1769),
    .VDD(VPWR),
    .Y(_03825_),
    .VSS(VGND),
    .A1(_03795_),
    .A2(_03823_));
 sg13g2_a21oi_1 _09710_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03795_),
    .A2(_03823_),
    .Y(_03826_),
    .B1(_03825_));
 sg13g2_nor2_1 _09711_ (.A(_03826_),
    .B(_03785_),
    .Y(_03827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _09712_ (.A(_03642_),
    .B_N(\acc_sum.add_renorm0.mantisa[10] ),
    .Y(_03828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1754 (.A(net1751),
    .X(net1754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09715_ (.A(\acc_sum.add_renorm0.exp[6] ),
    .B(net1690),
    .Y(_03831_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09716_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03831_),
    .Y(_03832_),
    .A2(_03820_),
    .A1(net1690));
 sg13g2_nand2_1 _09717_ (.Y(_03833_),
    .A(net1690),
    .B(_03796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09718_ (.B1(_03833_),
    .VDD(VPWR),
    .Y(_03834_),
    .VSS(VGND),
    .A1(_02924_),
    .A2(net1690));
 sg13g2_nor2_1 _09719_ (.A(\acc_sum.add_renorm0.exp[4] ),
    .B(net1690),
    .Y(_03835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09720_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03835_),
    .Y(_03836_),
    .A2(_03815_),
    .A1(net1690));
 sg13g2_nor2_1 _09721_ (.A(_03834_),
    .B(_03836_),
    .Y(_03837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09722_ (.Y(_03838_),
    .A(_03837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09723_ (.Y(_03839_),
    .A(_03828_),
    .B(\acc_sum.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09724_ (.Y(_03840_),
    .A(_02930_),
    .B(_03839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1698 (.A(_05046_),
    .X(net1698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09726_ (.Y(_03842_),
    .A(_03677_),
    .B(_03680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09727_ (.A(_03840_),
    .B(_03842_),
    .Y(_03843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09728_ (.Y(_03844_),
    .A(_02932_),
    .B(_03828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09729_ (.VDD(VPWR),
    .Y(_03845_),
    .A(_03844_),
    .VSS(VGND));
 sg13g2_xnor2_1 _09730_ (.Y(_03846_),
    .A(_03840_),
    .B(_03842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09731_ (.A(_03845_),
    .B(_03846_),
    .Y(_03847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09732_ (.Y(_03848_),
    .A(_03828_),
    .B(_03801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09733_ (.B1(_03848_),
    .VDD(VPWR),
    .Y(_03849_),
    .VSS(VGND),
    .A1(_02928_),
    .A2(_03828_));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09735_ (.Y(_03851_),
    .A(_03849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09736_ (.Y(_03852_),
    .A(_03851_),
    .B(_03678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09737_ (.B1(_03852_),
    .VDD(VPWR),
    .Y(_03853_),
    .VSS(VGND),
    .A1(_03843_),
    .A2(_03847_));
 sg13g2_nand2_1 _09738_ (.Y(_03854_),
    .A(_03678_),
    .B(_03849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _09739_ (.A(_03853_),
    .B(_03854_),
    .X(_03855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09740_ (.A(\acc_sum.add_renorm0.exp[3] ),
    .B(_03828_),
    .Y(_03856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _09741_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_03856_),
    .Y(_03857_),
    .A2(_03810_),
    .A1(_03828_));
 sg13g2_inv_2 _09742_ (.Y(_03858_),
    .A(_03857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09743_ (.Y(_03859_),
    .A(_03855_),
    .B(_03858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09744_ (.A(_03838_),
    .B(_03859_),
    .Y(_03860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09745_ (.VDD(VPWR),
    .Y(_03861_),
    .A(_03860_),
    .VSS(VGND));
 sg13g2_inv_1 _09746_ (.VDD(VPWR),
    .Y(_03862_),
    .A(_03793_),
    .VSS(VGND));
 sg13g2_nand2_1 _09747_ (.Y(_03863_),
    .A(_03862_),
    .B(net1690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09748_ (.B1(_03863_),
    .VDD(VPWR),
    .Y(_03864_),
    .VSS(VGND),
    .A1(_02920_),
    .A2(net1690));
 sg13g2_inv_2 _09749_ (.Y(_03865_),
    .A(_03864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09750_ (.B1(_03865_),
    .VDD(VPWR),
    .Y(_03866_),
    .VSS(VGND),
    .A1(_03832_),
    .A2(_03861_));
 sg13g2_inv_2 _09751_ (.Y(_03867_),
    .A(_03832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09752_ (.B(_03864_),
    .C(_03867_),
    .A(_03860_),
    .Y(_03868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09753_ (.B(net1664),
    .C(_03868_),
    .A(_03866_),
    .Y(_03869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09754_ (.Y(_03870_),
    .A(_03851_),
    .B(_03628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09755_ (.A(_03857_),
    .B(_03870_),
    .Y(_03871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09756_ (.VDD(VPWR),
    .Y(_03872_),
    .A(_03871_),
    .VSS(VGND));
 sg13g2_nor2_1 _09757_ (.A(_03838_),
    .B(_03872_),
    .Y(_03873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09758_ (.Y(_03874_),
    .A(_03873_),
    .B(_03867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09759_ (.Y(_03875_),
    .A(_03865_),
    .B(_03874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09760_ (.A(_03647_),
    .B(_03875_),
    .Y(_03876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09761_ (.VDD(VPWR),
    .Y(_03877_),
    .A(_03661_),
    .VSS(VGND));
 sg13g2_xnor2_1 _09762_ (.Y(_03878_),
    .A(_03851_),
    .B(_03661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09763_ (.A(_03840_),
    .B(_03878_),
    .Y(_03879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09764_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03877_),
    .A2(_03849_),
    .Y(_03880_),
    .B1(_03879_));
 sg13g2_nand2_1 _09765_ (.Y(_03881_),
    .A(_03880_),
    .B(_03858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09766_ (.A(_03838_),
    .B(_03881_),
    .Y(_03882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09767_ (.Y(_03883_),
    .A(_03882_),
    .B(_03867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09768_ (.B1(_03663_),
    .VDD(VPWR),
    .Y(_03884_),
    .VSS(VGND),
    .A1(_03865_),
    .A2(_03883_));
 sg13g2_a21oi_1 _09769_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03865_),
    .A2(_03883_),
    .Y(_03885_),
    .B1(_03884_));
 sg13g2_nor3_1 _09770_ (.A(net1769),
    .B(_03876_),
    .C(_03885_),
    .Y(_03886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09771_ (.Y(_03887_),
    .A(_03869_),
    .B(_03886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09772_ (.Y(_03888_),
    .A(_03827_),
    .B(_03887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09773_ (.Y(_03889_),
    .A(net1768),
    .B(\acc_sum.y[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09774_ (.Y(_01239_),
    .A(_03888_),
    .B(_03889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09775_ (.Y(_03890_),
    .A(_03861_),
    .B(_03867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09776_ (.Y(_03891_),
    .A(_03860_),
    .B(_03832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09777_ (.B(net1664),
    .C(_03891_),
    .A(_03890_),
    .Y(_03892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09778_ (.Y(_03893_),
    .A(_03867_),
    .B(_03873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09779_ (.Y(_03894_),
    .A(_03867_),
    .B(_03882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09780_ (.Y(_03895_),
    .B1(_03663_),
    .B2(_03894_),
    .A2(_03893_),
    .A1(_03648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09781_ (.B(_03895_),
    .C(net1803),
    .A(_03892_),
    .Y(_03896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09782_ (.A(_03822_),
    .B(_03819_),
    .Y(_03897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09783_ (.VDD(VPWR),
    .Y(_03898_),
    .A(_03823_),
    .VSS(VGND));
 sg13g2_o21ai_1 _09784_ (.B1(net1769),
    .VDD(VPWR),
    .Y(_03899_),
    .VSS(VGND),
    .A1(_03897_),
    .A2(_03898_));
 sg13g2_nand3_1 _09785_ (.B(_03783_),
    .C(_03899_),
    .A(_03896_),
    .Y(_03900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09786_ (.Y(_03901_),
    .A(_03782_),
    .B(\acc_sum.y[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09787_ (.Y(_01238_),
    .A(_03900_),
    .B(_03901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09788_ (.VDD(VPWR),
    .Y(_03902_),
    .A(_03819_),
    .VSS(VGND));
 sg13g2_nand2_1 _09789_ (.Y(_03903_),
    .A(_03818_),
    .B(_03799_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03902_),
    .A2(_03903_),
    .Y(_03904_),
    .B1(net1803));
 sg13g2_nand2b_1 _09791_ (.Y(_03905_),
    .B(_03783_),
    .A_N(_03904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09792_ (.VDD(VPWR),
    .Y(_03906_),
    .A(_03834_),
    .VSS(VGND));
 sg13g2_inv_1 _09793_ (.VDD(VPWR),
    .Y(_03907_),
    .A(_03881_),
    .VSS(VGND));
 sg13g2_inv_2 _09794_ (.Y(_03908_),
    .A(_03836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09795_ (.Y(_03909_),
    .A(_03907_),
    .B(_03908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09796_ (.VDD(VPWR),
    .Y(_03910_),
    .A(_03909_),
    .VSS(VGND));
 sg13g2_nor2_1 _09797_ (.A(_03906_),
    .B(_03910_),
    .Y(_03911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09798_ (.B1(_03663_),
    .VDD(VPWR),
    .Y(_03912_),
    .VSS(VGND),
    .A1(_03882_),
    .A2(_03911_));
 sg13g2_a21oi_1 _09799_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03871_),
    .A2(_03908_),
    .Y(_03913_),
    .B1(_03906_));
 sg13g2_o21ai_1 _09800_ (.B1(_03648_),
    .VDD(VPWR),
    .Y(_03914_),
    .VSS(VGND),
    .A1(_03873_),
    .A2(_03913_));
 sg13g2_nand3_1 _09801_ (.B(net1803),
    .C(_03914_),
    .A(_03912_),
    .Y(_03915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09802_ (.A(_03836_),
    .B(_03859_),
    .Y(_03916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09803_ (.A(_03906_),
    .B(_03916_),
    .Y(_03917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09804_ (.B1(net1664),
    .VDD(VPWR),
    .Y(_03918_),
    .VSS(VGND),
    .A1(_03860_),
    .A2(_03917_));
 sg13g2_nor2b_1 _09805_ (.A(_03915_),
    .B_N(_03918_),
    .Y(_03919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09806_ (.Y(_03920_),
    .A(net1768),
    .B(\acc_sum.y[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09807_ (.B1(_03920_),
    .VDD(VPWR),
    .Y(_01237_),
    .VSS(VGND),
    .A1(_03905_),
    .A2(_03919_));
 sg13g2_xnor2_1 _09808_ (.Y(_03921_),
    .A(_03836_),
    .B(_03871_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09809_ (.A(_03908_),
    .B(_03907_),
    .Y(_03922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09810_ (.B1(_03663_),
    .VDD(VPWR),
    .Y(_03923_),
    .VSS(VGND),
    .A1(_03922_),
    .A2(_03910_));
 sg13g2_o21ai_1 _09811_ (.B1(_03923_),
    .VDD(VPWR),
    .Y(_03924_),
    .VSS(VGND),
    .A1(_03647_),
    .A2(_03921_));
 sg13g2_inv_1 _09812_ (.VDD(VPWR),
    .Y(_03925_),
    .A(_03859_),
    .VSS(VGND));
 sg13g2_nor2_1 _09813_ (.A(_03908_),
    .B(_03925_),
    .Y(_03926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09814_ (.B1(net1664),
    .VDD(VPWR),
    .Y(_03927_),
    .VSS(VGND),
    .A1(_03916_),
    .A2(_03926_));
 sg13g2_nand3b_1 _09815_ (.B(_03927_),
    .C(net1803),
    .Y(_03928_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_03924_));
 sg13g2_nor2_1 _09816_ (.A(_03817_),
    .B(_03813_),
    .Y(_03929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09817_ (.VDD(VPWR),
    .Y(_03930_),
    .A(_03818_),
    .VSS(VGND));
 sg13g2_o21ai_1 _09818_ (.B1(net1769),
    .VDD(VPWR),
    .Y(_03931_),
    .VSS(VGND),
    .A1(_03929_),
    .A2(_03930_));
 sg13g2_nand3_1 _09819_ (.B(_03783_),
    .C(_03931_),
    .A(_03928_),
    .Y(_03932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09820_ (.Y(_03933_),
    .A(_03782_),
    .B(\acc_sum.y[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09821_ (.Y(_01236_),
    .A(_03932_),
    .B(_03933_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09822_ (.VDD(VPWR),
    .Y(_03934_),
    .A(\acc_sum.y[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09823_ (.A(_03858_),
    .B(_03855_),
    .Y(_03935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09824_ (.B1(net1664),
    .VDD(VPWR),
    .Y(_03936_),
    .VSS(VGND),
    .A1(_03935_),
    .A2(_03925_));
 sg13g2_a21oi_1 _09825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03851_),
    .A2(_03628_),
    .Y(_03937_),
    .B1(_03858_));
 sg13g2_o21ai_1 _09826_ (.B1(_03648_),
    .VDD(VPWR),
    .Y(_03938_),
    .VSS(VGND),
    .A1(_03871_),
    .A2(_03937_));
 sg13g2_nor2_1 _09827_ (.A(_03858_),
    .B(_03880_),
    .Y(_03939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09828_ (.B1(_03663_),
    .VDD(VPWR),
    .Y(_03940_),
    .VSS(VGND),
    .A1(_03939_),
    .A2(_03907_));
 sg13g2_nand4_1 _09829_ (.B(net1803),
    .C(_03938_),
    .A(_03936_),
    .Y(_03941_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03940_));
 sg13g2_nor2_1 _09830_ (.A(_03812_),
    .B(_03809_),
    .Y(_03942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09831_ (.B1(net1769),
    .VDD(VPWR),
    .Y(_03943_),
    .VSS(VGND),
    .A1(_03942_),
    .A2(_03813_));
 sg13g2_nand3_1 _09832_ (.B(_03783_),
    .C(_03943_),
    .A(_03941_),
    .Y(_03944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09833_ (.B1(_03944_),
    .VDD(VPWR),
    .Y(_01235_),
    .VSS(VGND),
    .A1(\acc_sum.reg3en.q[0] ),
    .A2(_03934_));
 sg13g2_inv_1 _09834_ (.VDD(VPWR),
    .Y(_03945_),
    .A(\acc_sum.y[9] ),
    .VSS(VGND));
 sg13g2_or3_1 _09835_ (.A(_03843_),
    .B(_03847_),
    .C(_03852_),
    .X(_03946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09836_ (.B(net1664),
    .C(_03853_),
    .A(_03946_),
    .Y(_03947_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09837_ (.A(_03628_),
    .B(_03851_),
    .Y(_03948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03684_),
    .A2(_03851_),
    .Y(_03949_),
    .B1(_03948_));
 sg13g2_nand2_1 _09839_ (.Y(_03950_),
    .A(_03878_),
    .B(_03840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _09840_ (.B(_03663_),
    .C(_03950_),
    .Y(_03951_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_03879_));
 sg13g2_nand4_1 _09841_ (.B(net1803),
    .C(_03949_),
    .A(_03947_),
    .Y(_03952_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03951_));
 sg13g2_and2_1 _09842_ (.A(_03808_),
    .B(_03804_),
    .X(_03953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09843_ (.B1(net1769),
    .VDD(VPWR),
    .Y(_03954_),
    .VSS(VGND),
    .A1(_03809_),
    .A2(_03953_));
 sg13g2_nand3_1 _09844_ (.B(_03952_),
    .C(_03954_),
    .A(_03783_),
    .Y(_03955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09845_ (.B1(_03955_),
    .VDD(VPWR),
    .Y(_01234_),
    .VSS(VGND),
    .A1(net1820),
    .A2(_03945_));
 sg13g2_inv_1 _09846_ (.VDD(VPWR),
    .Y(_03956_),
    .A(\acc_sum.y[8] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _09847_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03733_),
    .A2(_03806_),
    .Y(_03957_),
    .B1(_03805_));
 sg13g2_xnor2_1 _09848_ (.Y(_03958_),
    .A(\acc_sum.add_renorm0.exp[1] ),
    .B(_03957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09849_ (.A(_03840_),
    .B(_03648_),
    .Y(_03959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03662_),
    .A2(_03840_),
    .Y(_03960_),
    .B1(_03959_));
 sg13g2_nor2_1 _09851_ (.A(_03740_),
    .B(_03960_),
    .Y(_03961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09852_ (.Y(_03962_),
    .A(_03846_),
    .B(_03845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _09853_ (.B(net1664),
    .C(_03962_),
    .Y(_03963_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_03847_));
 sg13g2_a22oi_1 _09854_ (.Y(_03964_),
    .B1(_03961_),
    .B2(_03963_),
    .A2(_03958_),
    .A1(net1769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09855_ (.Y(_03965_),
    .A(_03783_),
    .B(_03964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09856_ (.B1(_03965_),
    .VDD(VPWR),
    .Y(_01233_),
    .VSS(VGND),
    .A1(net1820),
    .A2(_03956_));
 sg13g2_inv_1 _09857_ (.VDD(VPWR),
    .Y(_03966_),
    .A(\acc_sum.y[7] ),
    .VSS(VGND));
 sg13g2_xor2_1 _09858_ (.B(_03733_),
    .A(_03807_),
    .X(_03967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09859_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03665_),
    .A2(_03844_),
    .Y(_03968_),
    .B1(_03740_));
 sg13g2_nand2_1 _09860_ (.Y(_03969_),
    .A(net1664),
    .B(_03845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09861_ (.Y(_03970_),
    .B1(_03968_),
    .B2(_03969_),
    .A2(_03967_),
    .A1(net1769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09862_ (.Y(_03971_),
    .A(_03783_),
    .B(_03970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09863_ (.B1(_03971_),
    .VDD(VPWR),
    .Y(_01232_),
    .VSS(VGND),
    .A1(\acc_sum.reg3en.q[0] ),
    .A2(_03966_));
 sg13g2_nand2_1 _09864_ (.Y(_03972_),
    .A(net1768),
    .B(\acc_sum.y[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09865_ (.B1(_03972_),
    .VDD(VPWR),
    .Y(_01231_),
    .VSS(VGND),
    .A1(net1768),
    .A2(_03775_));
 sg13g2_nor2_1 _09866_ (.A(net1820),
    .B(\acc_sum.y[5] ),
    .Y(_03973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09867_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03722_),
    .A2(net1820),
    .Y(_01230_),
    .B1(_03973_));
 sg13g2_nand2_1 _09868_ (.Y(_03974_),
    .A(_03684_),
    .B(_03674_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09869_ (.Y(_03975_),
    .A(_03687_),
    .B(_03655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09870_ (.Y(_03976_),
    .A(_03649_),
    .B(_03652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09871_ (.Y(_03977_),
    .B1(_03631_),
    .B2(_03666_),
    .A2(_03635_),
    .A1(_03630_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _09872_ (.B(_03975_),
    .C(_03976_),
    .A(_03974_),
    .Y(_03978_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03977_));
 sg13g2_a21oi_1 _09873_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03978_),
    .A2(net1803),
    .Y(_03979_),
    .B1(_03743_));
 sg13g2_nor2_1 _09874_ (.A(net1820),
    .B(\acc_sum.y[4] ),
    .Y(_03980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09875_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03979_),
    .A2(net1820),
    .Y(_01229_),
    .B1(_03980_));
 sg13g2_mux2_1 _09876_ (.A0(\acc_sum.y[3] ),
    .A1(_03757_),
    .S(net1820),
    .X(_01228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _09877_ (.A0(\acc_sum.y[2] ),
    .A1(_03765_),
    .S(net1820),
    .X(_01227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09878_ (.Y(_03981_),
    .A(net1768),
    .B(\acc_sum.y[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09879_ (.B1(_03981_),
    .VDD(VPWR),
    .Y(_01226_),
    .VSS(VGND),
    .A1(net1768),
    .A2(_03779_));
 sg13g2_nand2_1 _09880_ (.Y(_03982_),
    .A(net1768),
    .B(\acc_sum.y[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09881_ (.B1(_03982_),
    .VDD(VPWR),
    .Y(_01225_),
    .VSS(VGND),
    .A1(net1768),
    .A2(_03747_));
 sg13g2_inv_2 _09882_ (.Y(_03983_),
    .A(\fp16_res_pipe.reg1en.d[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout52 (.A(net55),
    .X(net52),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _09884_ (.Y(_01224_),
    .B(net1767),
    .A_N(\fp16_res_pipe.reg_add_sub.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _09885_ (.A0(\fp16_res_pipe.op_sign_logic0.s_a ),
    .A1(\fp16_res_pipe.exp_mant_logic0.a[15] ),
    .S(net1831),
    .X(_01223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09886_ (.VDD(VPWR),
    .Y(_03985_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[15] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09887_ (.A(net1831),
    .B(\fp16_res_pipe.op_sign_logic0.s_b ),
    .Y(_03986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09888_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1831),
    .A2(_03985_),
    .Y(_01222_),
    .B1(_03986_));
 sg13g2_mux2_1 _09889_ (.A0(\fp16_res_pipe.op_sign_logic0.add_sub ),
    .A1(\fp16_res_pipe.reg_add_sub.q[0] ),
    .S(net1831),
    .X(_01221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09890_ (.VDD(VPWR),
    .Y(_03987_),
    .A(\fp16_res_pipe.seg_reg0.q[29] ),
    .VSS(VGND));
 sg13g2_inv_4 _09891_ (.A(\fp16_res_pipe.reg1en.q[0] ),
    .Y(_03988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout56 (.A(net71),
    .X(net56),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1772 (.A(net1771),
    .X(net1772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09894_ (.A(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .B(net1765),
    .Y(_03991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _09895_ (.Y(_03992_),
    .A(\fp16_res_pipe.exp_mant_logic0.a[14] ),
    .B(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09896_ (.VDD(VPWR),
    .Y(_03993_),
    .A(_03992_),
    .VSS(VGND));
 sg13g2_nor2_1 _09897_ (.A(\fp16_res_pipe.exp_mant_logic0.b[12] ),
    .B(_03593_),
    .Y(_03994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09898_ (.Y(_03995_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09899_ (.A(\fp16_res_pipe.exp_mant_logic0.a[12] ),
    .B(_03995_),
    .Y(_03996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09900_ (.A(_03994_),
    .B(_03996_),
    .Y(_03997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09901_ (.VDD(VPWR),
    .Y(_03998_),
    .A(_03997_),
    .VSS(VGND));
 sg13g2_nor2_1 _09902_ (.A(\fp16_res_pipe.exp_mant_logic0.b[13] ),
    .B(_03591_),
    .Y(_03999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09903_ (.VDD(VPWR),
    .Y(_04000_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[13] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09904_ (.A(\fp16_res_pipe.exp_mant_logic0.a[13] ),
    .B(_04000_),
    .Y(_04001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09905_ (.A(_03999_),
    .B(_04001_),
    .Y(_04002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09906_ (.VDD(VPWR),
    .Y(_04003_),
    .A(_04002_),
    .VSS(VGND));
 sg13g2_nor2_1 _09907_ (.A(\fp16_res_pipe.exp_mant_logic0.b[11] ),
    .B(_03595_),
    .Y(_04004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09908_ (.VDD(VPWR),
    .Y(_04005_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[11] ),
    .VSS(VGND));
 sg13g2_nor2_1 _09909_ (.A(\fp16_res_pipe.exp_mant_logic0.a[11] ),
    .B(_04005_),
    .Y(_04006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09910_ (.A(_04004_),
    .B(_04006_),
    .Y(_04007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09911_ (.VDD(VPWR),
    .Y(_04008_),
    .A(_04007_),
    .VSS(VGND));
 sg13g2_nor4_1 _09912_ (.A(_03993_),
    .B(_03998_),
    .C(_04003_),
    .D(_04008_),
    .Y(_04009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _09913_ (.B(\fp16_res_pipe.exp_mant_logic0.b[8] ),
    .A(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .X(_04010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09914_ (.VDD(VPWR),
    .Y(_04011_),
    .A(_04010_),
    .VSS(VGND));
 sg13g2_inv_2 _09915_ (.Y(_04012_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09916_ (.A(\fp16_res_pipe.exp_mant_logic0.a[7] ),
    .B(_04012_),
    .Y(_04013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09917_ (.Y(_04014_),
    .A(_04012_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09918_ (.VDD(VPWR),
    .Y(_04015_),
    .A(_04014_),
    .VSS(VGND));
 sg13g2_nor2_1 _09919_ (.A(_04013_),
    .B(_04015_),
    .Y(_04016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _09920_ (.Y(_04017_),
    .A(_04011_),
    .B(_04016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09921_ (.VDD(VPWR),
    .Y(_04018_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09922_ (.Y(_04019_),
    .A(_04018_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09923_ (.Y(_04020_),
    .A(_03597_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09924_ (.Y(_04021_),
    .A(_04019_),
    .B(_04020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09925_ (.VDD(VPWR),
    .Y(_04022_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09926_ (.Y(_04023_),
    .A(_04022_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _09927_ (.Y(_04024_),
    .A(_03599_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09928_ (.Y(_04025_),
    .A(_04023_),
    .B(_04024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09929_ (.A(_04021_),
    .B(_04025_),
    .Y(_04026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09930_ (.VDD(VPWR),
    .Y(_04027_),
    .A(_04026_),
    .VSS(VGND));
 sg13g2_nor2_1 _09931_ (.A(_04017_),
    .B(_04027_),
    .Y(_04028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09932_ (.Y(_04029_),
    .A(_04009_),
    .B(_04028_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout125 (.A(net127),
    .X(net125),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09934_ (.Y(_04031_),
    .A(net1703),
    .B(\fp16_res_pipe.exp_mant_logic0.a[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09935_ (.Y(_01220_),
    .B1(_03991_),
    .B2(_04031_),
    .A2(net1765),
    .A1(_03987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09936_ (.VDD(VPWR),
    .Y(_04032_),
    .A(\fp16_res_pipe.seg_reg0.q[28] ),
    .VSS(VGND));
 sg13g2_inv_1 _09937_ (.VDD(VPWR),
    .Y(_04033_),
    .A(_04020_),
    .VSS(VGND));
 sg13g2_inv_1 _09938_ (.VDD(VPWR),
    .Y(_04034_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _09939_ (.Y(_04035_),
    .A(_04034_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09940_ (.B1(_04035_),
    .VDD(VPWR),
    .Y(_04036_),
    .VSS(VGND),
    .A1(_04013_),
    .A2(_04010_));
 sg13g2_inv_1 _09941_ (.VDD(VPWR),
    .Y(_04037_),
    .A(_04023_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09942_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04036_),
    .A2(_04024_),
    .Y(_04038_),
    .B1(_04037_));
 sg13g2_o21ai_1 _09943_ (.B1(_04019_),
    .VDD(VPWR),
    .Y(_04039_),
    .VSS(VGND),
    .A1(_04033_),
    .A2(_04038_));
 sg13g2_nand2_1 _09944_ (.Y(_04040_),
    .A(_04039_),
    .B(_04009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _09945_ (.VDD(VPWR),
    .Y(_04041_),
    .A(_04004_),
    .VSS(VGND));
 sg13g2_inv_1 _09946_ (.VDD(VPWR),
    .Y(_04042_),
    .A(_03994_),
    .VSS(VGND));
 sg13g2_o21ai_1 _09947_ (.B1(_04042_),
    .VDD(VPWR),
    .Y(_04043_),
    .VSS(VGND),
    .A1(_03996_),
    .A2(_04041_));
 sg13g2_nor2_1 _09948_ (.A(_03993_),
    .B(_04003_),
    .Y(_04044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _09949_ (.A(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .B(_03589_),
    .Y(_04045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _09950_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_04044_),
    .C1(_04045_),
    .B1(_04043_),
    .A1(_03992_),
    .Y(_04046_),
    .A2(_03999_));
 sg13g2_nand2_2 _09951_ (.Y(_04047_),
    .A(_04040_),
    .B(_04046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _09952_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04047_),
    .A2(_03591_),
    .Y(_04048_),
    .B1(net1766));
 sg13g2_o21ai_1 _09953_ (.B1(_04048_),
    .VDD(VPWR),
    .Y(_04049_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.exp_mant_logic0.b[13] ),
    .A2(_04047_));
 sg13g2_o21ai_1 _09954_ (.B1(_04049_),
    .VDD(VPWR),
    .Y(_01219_),
    .VSS(VGND),
    .A1(_04032_),
    .A2(net1831));
 sg13g2_nand2_2 _09955_ (.Y(_04050_),
    .A(_04047_),
    .B(_04029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _09956_ (.Y(_04051_),
    .A(net1689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09957_ (.A(net1766),
    .B(_04051_),
    .Y(_04052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _09959_ (.A(_04052_),
    .Y(_04054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _09961_ (.A(net1766),
    .B(net1689),
    .Y(_04056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09964_ (.Y(_04059_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[12] ),
    .B2(net1682),
    .A2(net1766),
    .A1(\fp16_res_pipe.seg_reg0.q[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09965_ (.B1(_04059_),
    .VDD(VPWR),
    .Y(_01218_),
    .VSS(VGND),
    .A1(_03995_),
    .A2(_04054_));
 sg13g2_a22oi_1 _09966_ (.Y(_04060_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[11] ),
    .B2(_04056_),
    .A2(net1765),
    .A1(\fp16_res_pipe.seg_reg0.q[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09967_ (.B1(_04060_),
    .VDD(VPWR),
    .Y(_01217_),
    .VSS(VGND),
    .A1(_04005_),
    .A2(_04054_));
 sg13g2_a22oi_1 _09968_ (.Y(_04061_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[10] ),
    .B2(_04056_),
    .A2(net1765),
    .A1(\fp16_res_pipe.seg_reg0.q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09969_ (.B1(_04061_),
    .VDD(VPWR),
    .Y(_01216_),
    .VSS(VGND),
    .A1(_04018_),
    .A2(_04054_));
 sg13g2_nand2_1 _09970_ (.Y(_04062_),
    .A(_04052_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09971_ (.Y(_04063_),
    .A(_04056_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09972_ (.Y(_04064_),
    .A(net1765),
    .B(\fp16_res_pipe.seg_reg0.q[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09973_ (.B(_04063_),
    .C(_04064_),
    .A(_04062_),
    .Y(_01215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09974_ (.Y(_04065_),
    .A(_04052_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09975_ (.Y(_04066_),
    .A(_04056_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _09976_ (.Y(_04067_),
    .A(net1765),
    .B(\fp16_res_pipe.seg_reg0.q[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09977_ (.B(_04066_),
    .C(_04067_),
    .A(_04065_),
    .Y(_01214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _09978_ (.Y(_04068_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[7] ),
    .B2(_04056_),
    .A2(net1765),
    .A1(\fp16_res_pipe.seg_reg0.q[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09979_ (.B1(_04068_),
    .VDD(VPWR),
    .Y(_01213_),
    .VSS(VGND),
    .A1(_04012_),
    .A2(_04054_));
 sg13g2_nor4_1 _09980_ (.A(\fp16_res_pipe.exp_mant_logic0.a[10] ),
    .B(\fp16_res_pipe.exp_mant_logic0.a[9] ),
    .C(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .D(\fp16_res_pipe.exp_mant_logic0.a[7] ),
    .Y(_04069_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _09981_ (.A(\fp16_res_pipe.exp_mant_logic0.a[14] ),
    .B(\fp16_res_pipe.exp_mant_logic0.a[13] ),
    .C(\fp16_res_pipe.exp_mant_logic0.a[12] ),
    .D(\fp16_res_pipe.exp_mant_logic0.a[11] ),
    .Y(_04070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _09982_ (.A(\fp16_res_pipe.exp_mant_logic0.a[6] ),
    .B(\fp16_res_pipe.exp_mant_logic0.a[5] ),
    .C(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .D(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .Y(_04071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _09983_ (.A(\fp16_res_pipe.exp_mant_logic0.a[2] ),
    .B(\fp16_res_pipe.exp_mant_logic0.a[1] ),
    .C(\fp16_res_pipe.exp_mant_logic0.a[0] ),
    .Y(_04072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _09984_ (.B(_04070_),
    .C(_04071_),
    .A(_04069_),
    .Y(_04073_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04072_));
 sg13g2_buf_1 fanout67 (.A(net71),
    .X(net67),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _09986_ (.B(\fp16_res_pipe.reg1en.q[0] ),
    .C(_04073_),
    .A(_04047_),
    .Y(_04075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09987_ (.B1(_04075_),
    .VDD(VPWR),
    .Y(_01212_),
    .VSS(VGND),
    .A1(net1831),
    .A2(_03444_));
 sg13g2_inv_1 _09988_ (.VDD(VPWR),
    .Y(_04076_),
    .A(net1703),
    .VSS(VGND));
 sg13g2_a21oi_1 _09989_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04039_),
    .A2(_04007_),
    .Y(_04077_),
    .B1(_04004_));
 sg13g2_o21ai_1 _09990_ (.B1(_04042_),
    .VDD(VPWR),
    .Y(_04078_),
    .VSS(VGND),
    .A1(_03996_),
    .A2(_04077_));
 sg13g2_nand2_1 _09991_ (.Y(_04079_),
    .A(_04011_),
    .B(_04014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _09992_ (.B1(_04079_),
    .VDD(VPWR),
    .Y(_04080_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .A2(_04034_));
 sg13g2_inv_1 _09993_ (.VDD(VPWR),
    .Y(_04081_),
    .A(_04080_),
    .VSS(VGND));
 sg13g2_inv_1 _09994_ (.VDD(VPWR),
    .Y(_04082_),
    .A(_04024_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09995_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04082_),
    .A2(_04019_),
    .Y(_04083_),
    .B1(_04033_));
 sg13g2_o21ai_1 _09996_ (.B1(_04083_),
    .VDD(VPWR),
    .Y(_04084_),
    .VSS(VGND),
    .A1(_04027_),
    .A2(_04081_));
 sg13g2_a21oi_1 _09997_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04084_),
    .A2(_04007_),
    .Y(_04085_),
    .B1(_04006_));
 sg13g2_inv_1 _09998_ (.VDD(VPWR),
    .Y(_04086_),
    .A(_04085_),
    .VSS(VGND));
 sg13g2_a21oi_1 _09999_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04086_),
    .A2(_04042_),
    .Y(_04087_),
    .B1(_03996_));
 sg13g2_nor2_1 _10000_ (.A(_04051_),
    .B(_04087_),
    .Y(_04088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10001_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04078_),
    .A2(_04051_),
    .Y(_04089_),
    .B1(_04088_));
 sg13g2_xnor2_1 _10002_ (.Y(_04090_),
    .A(_04002_),
    .B(_04089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10003_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04078_),
    .A2(_04002_),
    .Y(_04091_),
    .B1(_03999_));
 sg13g2_nand2_1 _10004_ (.Y(_04092_),
    .A(_03589_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _10005_ (.B(_04092_),
    .C(_04029_),
    .Y(_04093_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_04091_));
 sg13g2_nor2_1 _10006_ (.A(_04003_),
    .B(_04087_),
    .Y(_04094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10007_ (.B1(_04050_),
    .VDD(VPWR),
    .Y(_04095_),
    .VSS(VGND),
    .A1(_04001_),
    .A2(_04094_));
 sg13g2_nand2_1 _10008_ (.Y(_04096_),
    .A(_04093_),
    .B(_04095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10009_ (.Y(_04097_),
    .A(_04096_),
    .B(_03993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10010_ (.Y(_04098_),
    .A(_04050_),
    .B(_04086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10011_ (.B1(_04098_),
    .VDD(VPWR),
    .Y(_04099_),
    .VSS(VGND),
    .A1(_04077_),
    .A2(_04050_));
 sg13g2_xnor2_1 _10012_ (.Y(_04100_),
    .A(_03998_),
    .B(_04099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _10013_ (.A0(_04039_),
    .A1(_04084_),
    .S(net1689),
    .X(_04101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10014_ (.Y(_04102_),
    .A(_04008_),
    .B(_04101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10015_ (.A(_04100_),
    .B(_04102_),
    .Y(_04103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10016_ (.Y(_04104_),
    .A(_04097_),
    .B(_04103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10017_ (.A(_04090_),
    .B(_04104_),
    .Y(_04105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_50_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_50_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10019_ (.Y(_04107_),
    .A(net1689),
    .B(_04014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10020_ (.B1(_04107_),
    .VDD(VPWR),
    .Y(_04108_),
    .VSS(VGND),
    .A1(_04013_),
    .A2(net1689));
 sg13g2_xnor2_1 _10021_ (.Y(_04109_),
    .A(_04010_),
    .B(_04108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10022_ (.A(_04016_),
    .B(_04109_),
    .Y(_04110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10023_ (.VDD(VPWR),
    .Y(_04111_),
    .A(_04110_),
    .VSS(VGND));
 sg13g2_nand2_1 _10024_ (.Y(_04112_),
    .A(net1689),
    .B(_04081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10025_ (.B1(_04112_),
    .VDD(VPWR),
    .Y(_04113_),
    .VSS(VGND),
    .A1(_04036_),
    .A2(net1689));
 sg13g2_xnor2_1 _10026_ (.Y(_04114_),
    .A(_04025_),
    .B(_04113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10027_ (.VDD(VPWR),
    .Y(_04115_),
    .A(_04114_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10028_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04081_),
    .A2(_04024_),
    .Y(_04116_),
    .B1(_04037_));
 sg13g2_nor2_1 _10029_ (.A(_04116_),
    .B(_04051_),
    .Y(_04117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04038_),
    .A2(_04051_),
    .Y(_04118_),
    .B1(_04117_));
 sg13g2_xor2_1 _10031_ (.B(_04118_),
    .A(_04021_),
    .X(_04119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10032_ (.VDD(VPWR),
    .Y(_04120_),
    .A(_04119_),
    .VSS(VGND));
 sg13g2_nor2_1 _10033_ (.A(_04115_),
    .B(_04120_),
    .Y(_04121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10034_ (.VDD(VPWR),
    .Y(_04122_),
    .A(_04121_),
    .VSS(VGND));
 sg13g2_nor2_1 _10035_ (.A(_04111_),
    .B(_04122_),
    .Y(_04123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10036_ (.Y(_04124_),
    .A(net1662),
    .B(_04123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_75_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_75_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10038_ (.Y(_04126_),
    .A(_04124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10039_ (.Y(_04127_),
    .B1(net1746),
    .B2(_04126_),
    .A2(net1688),
    .A1(net1827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10040_ (.A(_04114_),
    .B(_04120_),
    .Y(_04128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1876 (.A(net1875),
    .X(net1876),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10042_ (.Y(_04130_),
    .A(_04128_),
    .B(_04017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _10043_ (.B(_04097_),
    .C(_04103_),
    .Y(_04131_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_04090_));
 sg13g2_buf_8 clkbuf_leaf_47_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10045_ (.B1(net1703),
    .VDD(VPWR),
    .Y(_04133_),
    .VSS(VGND),
    .A1(_04130_),
    .A2(_04131_));
 sg13g2_nor3_1 _10046_ (.A(_04017_),
    .B(_04115_),
    .C(_04119_),
    .Y(_04134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10047_ (.Y(_04135_),
    .A(_04105_),
    .B(_04134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10048_ (.Y(_04136_),
    .A(_04124_),
    .B(_04135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10049_ (.VDD(VPWR),
    .Y(_04137_),
    .A(_04016_),
    .VSS(VGND));
 sg13g2_nand2_2 _10050_ (.Y(_04138_),
    .A(_04109_),
    .B(_04137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10051_ (.VDD(VPWR),
    .Y(_04139_),
    .A(_04138_),
    .VSS(VGND));
 sg13g2_nand3_1 _10052_ (.B(_04121_),
    .C(_04139_),
    .A(_04105_),
    .Y(_04140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_76_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_76_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10054_ (.A(_04011_),
    .B(_04137_),
    .Y(_04142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10055_ (.VDD(VPWR),
    .Y(_04143_),
    .A(_04142_),
    .VSS(VGND));
 sg13g2_nor2_1 _10056_ (.A(_04143_),
    .B(_04122_),
    .Y(_04144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10057_ (.VDD(VPWR),
    .Y(_04145_),
    .A(_04128_),
    .VSS(VGND));
 sg13g2_nor2_1 _10058_ (.A(_04017_),
    .B(_04145_),
    .Y(_04146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10059_ (.B1(_04105_),
    .VDD(VPWR),
    .Y(_04147_),
    .VSS(VGND),
    .A1(_04144_),
    .A2(_04146_));
 sg13g2_nand2_1 _10060_ (.Y(_04148_),
    .A(_04140_),
    .B(_04147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10061_ (.A(_04133_),
    .B(_04136_),
    .C(_04148_),
    .Y(_04149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10062_ (.A(_04054_),
    .B(_04149_),
    .Y(_04150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_99_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_99_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _10064_ (.Y(_04152_),
    .B(net1637),
    .A_N(_04127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout55 (.A(net56),
    .X(net55),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10066_ (.Y(_04154_),
    .B1(net1827),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[9] ),
    .A1(net1764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10067_ (.Y(_01211_),
    .A(_04152_),
    .B(_04154_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10068_ (.Y(_04155_),
    .A(_04126_),
    .B(net1827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10069_ (.Y(_04156_),
    .A(net1662),
    .B(_04144_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_77_clk (.A(clknet_5_27__leaf_clk),
    .X(clknet_leaf_77_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10071_ (.VDD(VPWR),
    .Y(_04158_),
    .A(_04156_),
    .VSS(VGND));
 sg13g2_nand2_1 _10072_ (.Y(_04159_),
    .A(net1643),
    .B(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10073_ (.Y(_04160_),
    .A(net1688),
    .B(net1828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10074_ (.B(_04159_),
    .C(_04160_),
    .A(_04155_),
    .Y(_04161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10075_ (.Y(_04162_),
    .A(net1637),
    .B(_04161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10076_ (.Y(_04163_),
    .B1(net1828),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[8] ),
    .A1(net1764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10077_ (.Y(_01210_),
    .A(_04162_),
    .B(_04163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10078_ (.Y(_04164_),
    .B1(net1827),
    .B2(net1643),
    .A2(net1688),
    .A1(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _10079_ (.A(_04140_),
    .Y(_04165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10080_ (.Y(_04166_),
    .A(_04165_),
    .B(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10081_ (.Y(_04167_),
    .A(_04126_),
    .B(net1828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10082_ (.B(_04166_),
    .C(_04167_),
    .A(_04164_),
    .Y(_04168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10083_ (.Y(_04169_),
    .A(_04168_),
    .B(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10084_ (.Y(_04170_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[7] ),
    .A1(net1764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10085_ (.Y(_01209_),
    .A(_04169_),
    .B(_04170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10086_ (.A(_03607_),
    .B(_04156_),
    .Y(_04171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10087_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .A2(_04126_),
    .Y(_04172_),
    .B1(_04171_));
 sg13g2_nand2_1 _10088_ (.Y(_04173_),
    .A(_04076_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10089_ (.Y(_04174_),
    .A(_04165_),
    .B(net1827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10090_ (.Y(_04175_),
    .A(net1662),
    .B(_04146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1670 (.A(_04530_),
    .X(net1670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _10092_ (.A(_04175_),
    .Y(_04177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10093_ (.Y(_04178_),
    .A(_04177_),
    .B(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _10094_ (.B(_04173_),
    .C(_04174_),
    .A(_04172_),
    .Y(_04179_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04178_));
 sg13g2_nand2_1 _10095_ (.Y(_04180_),
    .A(_04179_),
    .B(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10096_ (.Y(_04181_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[6] ),
    .A1(net1764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10097_ (.Y(_01208_),
    .A(_04180_),
    .B(_04181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10098_ (.A(_03613_),
    .B(net1703),
    .Y(_04182_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10099_ (.A(_03609_),
    .B(_04156_),
    .Y(_04183_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10100_ (.A(_03605_),
    .B(_04175_),
    .Y(_04184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10101_ (.A(_04182_),
    .B(_04183_),
    .C(_04184_),
    .Y(_04185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10102_ (.A(_03611_),
    .B(_04124_),
    .Y(_04186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10103_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04165_),
    .A2(net1828),
    .Y(_04187_),
    .B1(_04186_));
 sg13g2_nor2_1 _10104_ (.A(_04111_),
    .B(_04145_),
    .Y(_04188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10105_ (.Y(_04189_),
    .A(net1662),
    .B(_04188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10106_ (.Y(_04190_),
    .A(_04189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10107_ (.Y(_04191_),
    .A(net1642),
    .B(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10108_ (.B(_04187_),
    .C(_04191_),
    .A(_04185_),
    .Y(_04192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10109_ (.Y(_04193_),
    .A(_04192_),
    .B(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10110_ (.Y(_04194_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[2] ),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[5] ),
    .A1(net1764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10111_ (.Y(_01207_),
    .A(_04193_),
    .B(_04194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10112_ (.A(_04143_),
    .B(_04131_),
    .Y(_04195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10113_ (.B(net1746),
    .C(_04128_),
    .A(_04195_),
    .Y(_04196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10114_ (.B1(_04196_),
    .VDD(VPWR),
    .Y(_04197_),
    .VSS(VGND),
    .A1(_03611_),
    .A2(_04156_));
 sg13g2_nor2_1 _10115_ (.A(_03615_),
    .B(net1703),
    .Y(_04198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04177_),
    .A2(net1828),
    .Y(_04199_),
    .B1(_04198_));
 sg13g2_nor2b_1 _10117_ (.A(_04197_),
    .B_N(_04199_),
    .Y(_04200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10118_ (.A(_03605_),
    .B(_04189_),
    .Y(_04201_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10119_ (.A(_03613_),
    .B(_04124_),
    .Y(_04202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10120_ (.A(_03609_),
    .B(_04140_),
    .Y(_04203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10121_ (.A(_04201_),
    .B(_04202_),
    .C(_04203_),
    .Y(_04204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10122_ (.Y(_04205_),
    .A(_04200_),
    .B(_04204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10123_ (.Y(_04206_),
    .A(_04205_),
    .B(_04150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10124_ (.Y(_04207_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[1] ),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[4] ),
    .A1(net1763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10125_ (.Y(_01206_),
    .A(_04206_),
    .B(_04207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10126_ (.Y(_04208_),
    .A(net1642),
    .B(net1828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10127_ (.B1(_04208_),
    .VDD(VPWR),
    .Y(_04209_),
    .VSS(VGND),
    .A1(_03611_),
    .A2(_04140_));
 sg13g2_nor3_2 _10128_ (.A(_04145_),
    .B(_04138_),
    .C(_04131_),
    .Y(_04210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10129_ (.Y(_04211_),
    .A(_04210_),
    .B(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10130_ (.B1(_04211_),
    .VDD(VPWR),
    .Y(_04212_),
    .VSS(VGND),
    .A1(_03615_),
    .A2(_04124_));
 sg13g2_nor2_1 _10131_ (.A(_04209_),
    .B(_04212_),
    .Y(_04213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10132_ (.Y(_04214_),
    .A(net1643),
    .B(\fp16_res_pipe.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10133_ (.B1(_04214_),
    .VDD(VPWR),
    .Y(_04215_),
    .VSS(VGND),
    .A1(_03609_),
    .A2(_04175_));
 sg13g2_nand3_1 _10134_ (.B(net1827),
    .C(_04128_),
    .A(_04195_),
    .Y(_04216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10135_ (.B1(_04216_),
    .VDD(VPWR),
    .Y(_04217_),
    .VSS(VGND),
    .A1(_03617_),
    .A2(net1703));
 sg13g2_nor2_1 _10136_ (.A(_04215_),
    .B(_04217_),
    .Y(_04218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10137_ (.Y(_04219_),
    .A(_04213_),
    .B(_04218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10138_ (.Y(_04220_),
    .A(_04219_),
    .B(_04150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10139_ (.Y(_04221_),
    .B1(\fp16_res_pipe.exp_mant_logic0.a[0] ),
    .B2(net1682),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_a[3] ),
    .A1(net1763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10140_ (.Y(_01205_),
    .A(_04220_),
    .B(_04221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10141_ (.B(_04128_),
    .C(_04139_),
    .A(net1662),
    .Y(_04222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_78_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_78_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10143_ (.Y(_04224_),
    .A(_04135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10144_ (.Y(_04225_),
    .A(_04224_),
    .B(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10145_ (.B1(_04225_),
    .VDD(VPWR),
    .Y(_04226_),
    .VSS(VGND),
    .A1(_03605_),
    .A2(_04222_));
 sg13g2_nand3_1 _10146_ (.B(_04128_),
    .C(_04142_),
    .A(net1662),
    .Y(_04227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_79_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_79_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10148_ (.Y(_04229_),
    .A(net1642),
    .B(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10149_ (.B1(_04229_),
    .VDD(VPWR),
    .Y(_04230_),
    .VSS(VGND),
    .A1(_03607_),
    .A2(_04227_));
 sg13g2_nor2_1 _10150_ (.A(_04226_),
    .B(_04230_),
    .Y(_04231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10151_ (.A(_04138_),
    .B(_04122_),
    .Y(_04232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10152_ (.Y(_04233_),
    .A(net1662),
    .B(_04232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_80_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_80_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10154_ (.Y(_04235_),
    .A(_04177_),
    .B(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10155_ (.B1(_04235_),
    .VDD(VPWR),
    .Y(_04236_),
    .VSS(VGND),
    .A1(_03613_),
    .A2(_04233_));
 sg13g2_nand2_1 _10156_ (.Y(_04237_),
    .A(net1643),
    .B(\fp16_res_pipe.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10157_ (.B1(_04237_),
    .VDD(VPWR),
    .Y(_04238_),
    .VSS(VGND),
    .A1(_03617_),
    .A2(_04124_));
 sg13g2_nor2_1 _10158_ (.A(_04236_),
    .B(_04238_),
    .Y(_04239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10159_ (.Y(_04240_),
    .A(_04231_),
    .B(_04239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10160_ (.Y(_04241_),
    .A(_04240_),
    .B(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10161_ (.Y(_04242_),
    .A(net1764),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10162_ (.Y(_01204_),
    .A(_04241_),
    .B(_04242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10163_ (.Y(_04243_),
    .A(_04224_),
    .B(net1827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10164_ (.B1(_04243_),
    .VDD(VPWR),
    .Y(_04244_),
    .VSS(VGND),
    .A1(_03607_),
    .A2(_04222_));
 sg13g2_nand2_1 _10165_ (.Y(_04245_),
    .A(net1642),
    .B(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10166_ (.B1(_04245_),
    .VDD(VPWR),
    .Y(_04246_),
    .VSS(VGND),
    .A1(_03609_),
    .A2(_04227_));
 sg13g2_nor2_1 _10167_ (.A(_04244_),
    .B(_04246_),
    .Y(_04247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10168_ (.A(_03613_),
    .B(_04175_),
    .Y(_04248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10169_ (.A(_03617_),
    .B(_04156_),
    .Y(_04249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10170_ (.A(_03615_),
    .B(_04233_),
    .Y(_04250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10171_ (.A(_04248_),
    .B(_04249_),
    .C(_04250_),
    .Y(_04251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10172_ (.Y(_04252_),
    .A(_04247_),
    .B(_04251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10173_ (.Y(_04253_),
    .A(_04252_),
    .B(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10174_ (.Y(_04254_),
    .A(net1764),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10175_ (.Y(_01203_),
    .A(_04253_),
    .B(_04254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10176_ (.A(_03611_),
    .B(_04227_),
    .Y(_04255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10177_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fp16_res_pipe.exp_mant_logic0.a[2] ),
    .A2(net1642),
    .Y(_04256_),
    .B1(_04255_));
 sg13g2_nor2_1 _10178_ (.A(_03609_),
    .B(_04222_),
    .Y(_04257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10179_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1828),
    .A2(_04224_),
    .Y(_04258_),
    .B1(_04257_));
 sg13g2_nor2_1 _10180_ (.A(_03617_),
    .B(_04233_),
    .Y(_04259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fp16_res_pipe.exp_mant_logic0.a[1] ),
    .A2(_04177_),
    .Y(_04260_),
    .B1(_04259_));
 sg13g2_nand3_1 _10182_ (.B(_04258_),
    .C(_04260_),
    .A(_04256_),
    .Y(_04261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10183_ (.Y(_04262_),
    .A(_04261_),
    .B(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10184_ (.Y(_04263_),
    .A(net1764),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10185_ (.Y(_01202_),
    .A(_04262_),
    .B(_04263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _10186_ (.A(\fp16_res_pipe.exp_mant_logic0.b[10] ),
    .B(\fp16_res_pipe.exp_mant_logic0.b[9] ),
    .C(\fp16_res_pipe.exp_mant_logic0.b[8] ),
    .D(\fp16_res_pipe.exp_mant_logic0.b[7] ),
    .Y(_04264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _10187_ (.A(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .B(\fp16_res_pipe.exp_mant_logic0.b[13] ),
    .C(\fp16_res_pipe.exp_mant_logic0.b[12] ),
    .D(\fp16_res_pipe.exp_mant_logic0.b[11] ),
    .Y(_04265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _10188_ (.A(\fp16_res_pipe.exp_mant_logic0.b[6] ),
    .B(\fp16_res_pipe.exp_mant_logic0.b[5] ),
    .C(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .D(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .Y(_04266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10189_ (.A(\fp16_res_pipe.exp_mant_logic0.b[2] ),
    .B(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .C(\fp16_res_pipe.exp_mant_logic0.b[0] ),
    .Y(_04267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _10190_ (.B(_04265_),
    .C(_04266_),
    .A(_04264_),
    .Y(_04268_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04267_));
 sg13g2_buf_2 fanout68 (.A(net70),
    .X(net68),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10192_ (.B(net1831),
    .C(_04268_),
    .A(net1689),
    .Y(_04270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10193_ (.B1(_04270_),
    .VDD(VPWR),
    .Y(_01201_),
    .VSS(VGND),
    .A1(net1831),
    .A2(_03368_));
 sg13g2_a22oi_1 _10194_ (.Y(_04271_),
    .B1(net1745),
    .B2(net1644),
    .A2(net1688),
    .A1(net1829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _10195_ (.A(_04149_),
    .B_N(_04056_),
    .Y(_04272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_100_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_100_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _10197_ (.Y(_04274_),
    .B(net1636),
    .A_N(_04271_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10198_ (.Y(_04275_),
    .B1(net1829),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[9] ),
    .A1(_03988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10199_ (.Y(_01200_),
    .A(_04274_),
    .B(_04275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10200_ (.Y(_04276_),
    .A(net1644),
    .B(net1829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10201_ (.Y(_04277_),
    .A(net1643),
    .B(net1745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10202_ (.Y(_04278_),
    .A(net1688),
    .B(net1830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10203_ (.B(_04277_),
    .C(_04278_),
    .A(_04276_),
    .Y(_04279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10204_ (.Y(_04280_),
    .A(net1636),
    .B(_04279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10205_ (.Y(_04281_),
    .B1(net1830),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[8] ),
    .A1(_03988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10206_ (.Y(_01199_),
    .A(_04280_),
    .B(_04281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10207_ (.Y(_04282_),
    .B1(net1829),
    .B2(net1643),
    .A2(net1688),
    .A1(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10208_ (.Y(_04283_),
    .A(_04165_),
    .B(net1745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10209_ (.Y(_04284_),
    .A(net1644),
    .B(net1830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10210_ (.B(_04283_),
    .C(_04284_),
    .A(_04282_),
    .Y(_04285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10211_ (.Y(_04286_),
    .A(_04285_),
    .B(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10212_ (.Y(_04287_),
    .B1(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[7] ),
    .A1(net1763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10213_ (.Y(_01198_),
    .A(_04286_),
    .B(_04287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10214_ (.Y(_04288_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10215_ (.A(_04288_),
    .B(_04156_),
    .Y(_04289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .A2(net1644),
    .Y(_04290_),
    .B1(_04289_));
 sg13g2_nand2_1 _10217_ (.Y(_04291_),
    .A(net1688),
    .B(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10218_ (.Y(_04292_),
    .A(_04165_),
    .B(net1829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10219_ (.Y(_04293_),
    .A(_04177_),
    .B(net1745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _10220_ (.B(_04291_),
    .C(_04292_),
    .A(_04290_),
    .Y(_04294_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04293_));
 sg13g2_nand2_1 _10221_ (.Y(_04295_),
    .A(_04294_),
    .B(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10222_ (.Y(_04296_),
    .B1(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[6] ),
    .A1(net1763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10223_ (.Y(_01197_),
    .A(_04295_),
    .B(_04296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10224_ (.Y(_04297_),
    .B1(_04190_),
    .B2(net1745),
    .A2(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .A1(net1644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _10225_ (.A(\fp16_res_pipe.exp_mant_logic0.b[2] ),
    .Y(_04298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10226_ (.A(_04298_),
    .B(net1703),
    .Y(_04299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10227_ (.Y(_04300_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10228_ (.A(_04300_),
    .B(_04156_),
    .Y(_04301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10229_ (.Y(_04302_),
    .A(net1829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10230_ (.A(_04302_),
    .B(_04175_),
    .Y(_04303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10231_ (.A(_04299_),
    .B(_04301_),
    .C(_04303_),
    .Y(_04304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10232_ (.Y(_04305_),
    .A(_04165_),
    .B(net1830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10233_ (.B(_04304_),
    .C(_04305_),
    .A(_04297_),
    .Y(_04306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10234_ (.Y(_04307_),
    .A(_04306_),
    .B(_04272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10235_ (.Y(_04308_),
    .B1(\fp16_res_pipe.exp_mant_logic0.b[2] ),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[5] ),
    .A1(_03988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10236_ (.Y(_01196_),
    .A(_04307_),
    .B(_04308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10237_ (.A(_04302_),
    .B(_04189_),
    .Y(_04309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10238_ (.A(_04298_),
    .B(_04124_),
    .Y(_04310_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10239_ (.A(_04300_),
    .B(_04140_),
    .Y(_04311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10240_ (.A(_04309_),
    .B(_04310_),
    .C(_04311_),
    .Y(_04312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10241_ (.B(_04128_),
    .C(net1745),
    .A(_04195_),
    .Y(_04313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10242_ (.Y(_04314_),
    .A(net1688),
    .B(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10243_ (.A(_04313_),
    .B(_04314_),
    .X(_04315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10244_ (.Y(_04316_),
    .B1(net1830),
    .B2(_04177_),
    .A2(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .A1(net1643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10245_ (.B(_04315_),
    .C(_04316_),
    .A(_04312_),
    .Y(_04317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10246_ (.Y(_04318_),
    .A(_04317_),
    .B(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10247_ (.Y(_04319_),
    .B1(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[4] ),
    .A1(_03988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10248_ (.Y(_01195_),
    .A(_04318_),
    .B(_04319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10249_ (.Y(_04320_),
    .A(_04158_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10250_ (.B1(_04320_),
    .VDD(VPWR),
    .Y(_04321_),
    .VSS(VGND),
    .A1(_04300_),
    .A2(_04175_));
 sg13g2_inv_2 _10251_ (.Y(_04322_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10252_ (.B(net1829),
    .C(_04128_),
    .A(_04195_),
    .Y(_04323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10253_ (.B1(_04323_),
    .VDD(VPWR),
    .Y(_04324_),
    .VSS(VGND),
    .A1(_04322_),
    .A2(net1703));
 sg13g2_nor2_1 _10254_ (.A(_04321_),
    .B(_04324_),
    .Y(_04325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10255_ (.Y(_04326_),
    .A(_04210_),
    .B(net1745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10256_ (.Y(_04327_),
    .A(_04190_),
    .B(net1830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10257_ (.Y(_04328_),
    .A(_04326_),
    .B(_04327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10258_ (.Y(_04329_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10259_ (.Y(_04330_),
    .A(net1644),
    .B(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10260_ (.B1(_04330_),
    .VDD(VPWR),
    .Y(_04331_),
    .VSS(VGND),
    .A1(_04329_),
    .A2(_04140_));
 sg13g2_nor2_1 _10261_ (.A(_04328_),
    .B(_04331_),
    .Y(_04332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10262_ (.Y(_04333_),
    .A(_04325_),
    .B(_04332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10263_ (.Y(_04334_),
    .A(_04333_),
    .B(_04272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10264_ (.Y(_04335_),
    .B1(\fp16_res_pipe.exp_mant_logic0.b[0] ),
    .B2(net1683),
    .A2(\fp16_res_pipe.op_sign_logic0.mantisa_b[3] ),
    .A1(_03988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10265_ (.Y(_01194_),
    .A(_04334_),
    .B(_04335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10266_ (.Y(_04336_),
    .A(_04224_),
    .B(net1745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10267_ (.B1(_04336_),
    .VDD(VPWR),
    .Y(_04337_),
    .VSS(VGND),
    .A1(_04302_),
    .A2(_04222_));
 sg13g2_nand2_1 _10268_ (.Y(_04338_),
    .A(_04190_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10269_ (.B1(_04338_),
    .VDD(VPWR),
    .Y(_04339_),
    .VSS(VGND),
    .A1(_04288_),
    .A2(_04227_));
 sg13g2_nor2_1 _10270_ (.A(_04337_),
    .B(_04339_),
    .Y(_04340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10271_ (.Y(_04341_),
    .A(_04177_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10272_ (.B1(_04341_),
    .VDD(VPWR),
    .Y(_04342_),
    .VSS(VGND),
    .A1(_04298_),
    .A2(_04233_));
 sg13g2_nand2_1 _10273_ (.Y(_04343_),
    .A(net1643),
    .B(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10274_ (.B1(_04343_),
    .VDD(VPWR),
    .Y(_04344_),
    .VSS(VGND),
    .A1(_04322_),
    .A2(_04124_));
 sg13g2_nor2_1 _10275_ (.A(_04342_),
    .B(_04344_),
    .Y(_04345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10276_ (.Y(_04346_),
    .A(_04340_),
    .B(_04345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10277_ (.Y(_04347_),
    .A(_04346_),
    .B(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10278_ (.Y(_04348_),
    .A(net1763),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10279_ (.Y(_01193_),
    .A(_04347_),
    .B(_04348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10280_ (.Y(_04349_),
    .A(_04190_),
    .B(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10281_ (.B1(_04349_),
    .VDD(VPWR),
    .Y(_04350_),
    .VSS(VGND),
    .A1(_04300_),
    .A2(_04227_));
 sg13g2_a22oi_1 _10282_ (.Y(_04351_),
    .B1(net1830),
    .B2(_04210_),
    .A2(_04224_),
    .A1(net1829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10283_ (.A(_04322_),
    .B(_04156_),
    .Y(_04352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10284_ (.A(_04298_),
    .B(_04175_),
    .Y(_04353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10285_ (.VDD(VPWR),
    .Y(_04354_),
    .A(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10286_ (.A(_04354_),
    .B(_04233_),
    .Y(_04355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10287_ (.A(_04352_),
    .B(_04353_),
    .C(_04355_),
    .Y(_04356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _10288_ (.B(_04351_),
    .C(_04356_),
    .Y(_04357_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_04350_));
 sg13g2_nand2_1 _10289_ (.Y(_04358_),
    .A(_04357_),
    .B(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10290_ (.Y(_04359_),
    .A(net1763),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10291_ (.Y(_01192_),
    .A(_04358_),
    .B(_04359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10292_ (.Y(_04360_),
    .B1(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .B2(_04210_),
    .A2(_04224_),
    .A1(net1830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10293_ (.A(_04298_),
    .B(_04189_),
    .Y(_04361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10294_ (.A(_04329_),
    .B(_04227_),
    .Y(_04362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10295_ (.A(_04361_),
    .B(_04362_),
    .Y(_04363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10296_ (.A(_04322_),
    .B(_04233_),
    .Y(_04364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10297_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .A2(_04177_),
    .Y(_04365_),
    .B1(_04364_));
 sg13g2_nand3_1 _10298_ (.B(_04363_),
    .C(_04365_),
    .A(_04360_),
    .Y(_04366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10299_ (.Y(_04367_),
    .A(_04366_),
    .B(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10300_ (.Y(_04368_),
    .A(net1763),
    .B(\fp16_res_pipe.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10301_ (.Y(_01191_),
    .A(_04367_),
    .B(_04368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10302_ (.Y(_04369_),
    .A(net1911),
    .B(\fp16_res_pipe.x2[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10303_ (.B1(_04369_),
    .VDD(VPWR),
    .Y(_01190_),
    .VSS(VGND),
    .A1(net1911),
    .A2(_03985_));
 sg13g2_mux2_1 _10304_ (.A0(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .A1(\fp16_res_pipe.x2[14] ),
    .S(net1913),
    .X(_01189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10305_ (.Y(_04370_),
    .A(net1912),
    .B(\fp16_res_pipe.x2[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10306_ (.B1(_04370_),
    .VDD(VPWR),
    .Y(_01188_),
    .VSS(VGND),
    .A1(net1915),
    .A2(_04000_));
 sg13g2_nand2_1 _10307_ (.Y(_04371_),
    .A(net1914),
    .B(\fp16_res_pipe.x2[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10308_ (.B1(_04371_),
    .VDD(VPWR),
    .Y(_01187_),
    .VSS(VGND),
    .A1(net1915),
    .A2(_03995_));
 sg13g2_nand2_1 _10309_ (.Y(_04372_),
    .A(net1914),
    .B(\fp16_res_pipe.x2[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10310_ (.B1(_04372_),
    .VDD(VPWR),
    .Y(_01186_),
    .VSS(VGND),
    .A1(net1914),
    .A2(_04005_));
 sg13g2_nand2_1 _10311_ (.Y(_04373_),
    .A(net1912),
    .B(\fp16_res_pipe.x2[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10312_ (.B1(_04373_),
    .VDD(VPWR),
    .Y(_01185_),
    .VSS(VGND),
    .A1(net1914),
    .A2(_04018_));
 sg13g2_nand2_1 _10313_ (.Y(_04374_),
    .A(net1920),
    .B(\fp16_res_pipe.x2[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10314_ (.B1(_04374_),
    .VDD(VPWR),
    .Y(_01184_),
    .VSS(VGND),
    .A1(net1919),
    .A2(_04022_));
 sg13g2_nand2_1 _10315_ (.Y(_04375_),
    .A(net1912),
    .B(\fp16_res_pipe.x2[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10316_ (.B1(_04375_),
    .VDD(VPWR),
    .Y(_01183_),
    .VSS(VGND),
    .A1(net1919),
    .A2(_04034_));
 sg13g2_nand2_1 _10317_ (.Y(_04376_),
    .A(net1911),
    .B(\fp16_res_pipe.x2[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10318_ (.B1(_04376_),
    .VDD(VPWR),
    .Y(_01182_),
    .VSS(VGND),
    .A1(net1919),
    .A2(_04012_));
 sg13g2_nand2_1 _10319_ (.Y(_04377_),
    .A(net1920),
    .B(\fp16_res_pipe.x2[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10320_ (.B1(_04377_),
    .VDD(VPWR),
    .Y(_01181_),
    .VSS(VGND),
    .A1(net1919),
    .A2(_04302_));
 sg13g2_nand2_1 _10321_ (.Y(_04378_),
    .A(net1921),
    .B(\fp16_res_pipe.x2[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10322_ (.B1(_04378_),
    .VDD(VPWR),
    .Y(_01180_),
    .VSS(VGND),
    .A1(net1921),
    .A2(_04288_));
 sg13g2_nand2_1 _10323_ (.Y(_04379_),
    .A(net1920),
    .B(\fp16_res_pipe.x2[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10324_ (.B1(_04379_),
    .VDD(VPWR),
    .Y(_01179_),
    .VSS(VGND),
    .A1(net1921),
    .A2(_04300_));
 sg13g2_nand2_1 _10325_ (.Y(_04380_),
    .A(net1920),
    .B(\fp16_res_pipe.x2[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10326_ (.B1(_04380_),
    .VDD(VPWR),
    .Y(_01178_),
    .VSS(VGND),
    .A1(net1921),
    .A2(_04329_));
 sg13g2_nand2_1 _10327_ (.Y(_04381_),
    .A(net1921),
    .B(\fp16_res_pipe.x2[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10328_ (.B1(_04381_),
    .VDD(VPWR),
    .Y(_01177_),
    .VSS(VGND),
    .A1(net1921),
    .A2(_04298_));
 sg13g2_nand2_1 _10329_ (.Y(_04382_),
    .A(net1920),
    .B(\fp16_res_pipe.x2[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10330_ (.B1(_04382_),
    .VDD(VPWR),
    .Y(_01176_),
    .VSS(VGND),
    .A1(net1915),
    .A2(_04354_));
 sg13g2_nand2_1 _10331_ (.Y(_04383_),
    .A(net1921),
    .B(\fp16_res_pipe.x2[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10332_ (.B1(_04383_),
    .VDD(VPWR),
    .Y(_01175_),
    .VSS(VGND),
    .A1(net1921),
    .A2(_04322_));
 sg13g2_xor2_1 _10333_ (.B(\fp16_sum_pipe.op_sign_logic0.s_b ),
    .A(\fp16_sum_pipe.op_sign_logic0.s_a ),
    .X(_04384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1824 (.A(net1823),
    .X(net1824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10335_ (.Y(_04386_),
    .A(_04384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout84 (.A(net85),
    .X(net84),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10337_ (.A(\fp16_sum_pipe.seg_reg1.q[21] ),
    .B(net1844),
    .Y(_04388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10338_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04386_),
    .A2(net1844),
    .Y(_01174_),
    .B1(_04388_));
 sg13g2_inv_1 _10339_ (.VDD(VPWR),
    .Y(_04389_),
    .A(\fp16_sum_pipe.seg_reg1.q[20] ),
    .VSS(VGND));
 sg13g2_inv_1 _10340_ (.VDD(VPWR),
    .Y(_04390_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10341_ (.Y(_04391_),
    .A(_04390_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10342_ (.VDD(VPWR),
    .Y(_04392_),
    .A(_04391_),
    .VSS(VGND));
 sg13g2_inv_1 _10343_ (.VDD(VPWR),
    .Y(_04393_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[9] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10344_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[9] ),
    .B(_04393_),
    .Y(_04394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10345_ (.Y(_04395_),
    .A(_04393_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10346_ (.VDD(VPWR),
    .Y(_04396_),
    .A(_04395_),
    .VSS(VGND));
 sg13g2_nor2_2 _10347_ (.A(_04394_),
    .B(_04396_),
    .Y(_04397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10348_ (.VDD(VPWR),
    .Y(_04398_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[7] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10349_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[7] ),
    .B(_04398_),
    .Y(_04399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10350_ (.Y(_04400_),
    .A(_04398_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10351_ (.VDD(VPWR),
    .Y(_04401_),
    .A(_04400_),
    .VSS(VGND));
 sg13g2_nor2_1 _10352_ (.A(_04399_),
    .B(_04401_),
    .Y(_04402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10353_ (.Y(_04403_),
    .A(_04402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10354_ (.VDD(VPWR),
    .Y(_04404_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[6] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10355_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[6] ),
    .B(_04404_),
    .Y(_04405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10356_ (.Y(_04406_),
    .A(_04404_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10357_ (.Y(_04407_),
    .A(_04406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10358_ (.A(_04405_),
    .B(_04407_),
    .Y(_04408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10359_ (.VDD(VPWR),
    .Y(_04409_),
    .A(_04408_),
    .VSS(VGND));
 sg13g2_nor2_1 _10360_ (.A(_04403_),
    .B(_04409_),
    .Y(_04410_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10361_ (.VDD(VPWR),
    .Y(_04411_),
    .A(_04410_),
    .VSS(VGND));
 sg13g2_nand2b_2 _10362_ (.Y(_04412_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\fp16_sum_pipe.op_sign_logic0.mantisa_b[1] ));
 sg13g2_inv_1 _10363_ (.VDD(VPWR),
    .Y(_04413_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10364_ (.Y(_04414_),
    .A(_04413_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10365_ (.VDD(VPWR),
    .Y(_04415_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10366_ (.Y(_04416_),
    .A(_04415_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10367_ (.VDD(VPWR),
    .Y(_04417_),
    .A(_04416_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10368_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04412_),
    .A2(_04414_),
    .Y(_04418_),
    .B1(_04417_));
 sg13g2_inv_1 _10369_ (.VDD(VPWR),
    .Y(_04419_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[2] ),
    .VSS(VGND));
 sg13g2_nor2_2 _10370_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[2] ),
    .B(_04419_),
    .Y(_04420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10371_ (.Y(_04421_),
    .A(_04419_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10372_ (.VDD(VPWR),
    .Y(_04422_),
    .A(_04421_),
    .VSS(VGND));
 sg13g2_nor2_2 _10373_ (.A(_04420_),
    .B(_04422_),
    .Y(_04423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10374_ (.VDD(VPWR),
    .Y(_04424_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10375_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[3] ),
    .B(_04424_),
    .Y(_04425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10376_ (.Y(_04426_),
    .A(_04424_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10377_ (.VDD(VPWR),
    .Y(_04427_),
    .A(_04426_),
    .VSS(VGND));
 sg13g2_nor2_2 _10378_ (.A(_04425_),
    .B(_04427_),
    .Y(_04428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10379_ (.Y(_04429_),
    .A(_04423_),
    .B(_04428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10380_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04428_),
    .A2(_04420_),
    .Y(_04430_),
    .B1(_04427_));
 sg13g2_o21ai_1 _10381_ (.B1(_04430_),
    .VDD(VPWR),
    .Y(_04431_),
    .VSS(VGND),
    .A1(_04418_),
    .A2(_04429_));
 sg13g2_inv_1 _10382_ (.VDD(VPWR),
    .Y(_04432_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[4] ),
    .VSS(VGND));
 sg13g2_nor2_2 _10383_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[4] ),
    .B(_04432_),
    .Y(_04433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10384_ (.Y(_04434_),
    .A(_04432_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10385_ (.VDD(VPWR),
    .Y(_04435_),
    .A(_04434_),
    .VSS(VGND));
 sg13g2_nor2_2 _10386_ (.A(_04433_),
    .B(_04435_),
    .Y(_04436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10387_ (.VDD(VPWR),
    .Y(_04437_),
    .A(_04436_),
    .VSS(VGND));
 sg13g2_inv_1 _10388_ (.VDD(VPWR),
    .Y(_04438_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[5] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10389_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[5] ),
    .B(_04438_),
    .Y(_04439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10390_ (.Y(_04440_),
    .A(_04438_),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10391_ (.VDD(VPWR),
    .Y(_04441_),
    .A(_04440_),
    .VSS(VGND));
 sg13g2_nor2_1 _10392_ (.A(_04439_),
    .B(_04441_),
    .Y(_04442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10393_ (.VDD(VPWR),
    .Y(_04443_),
    .A(_04442_),
    .VSS(VGND));
 sg13g2_nor2_1 _10394_ (.A(_04437_),
    .B(_04443_),
    .Y(_04444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10395_ (.Y(_04445_),
    .A(_04431_),
    .B(_04444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10396_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04442_),
    .A2(_04433_),
    .Y(_04446_),
    .B1(_04441_));
 sg13g2_nand2_1 _10397_ (.Y(_04447_),
    .A(_04445_),
    .B(_04446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10398_ (.VDD(VPWR),
    .Y(_04448_),
    .A(_04447_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10399_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04402_),
    .A2(_04407_),
    .Y(_04449_),
    .B1(_04401_));
 sg13g2_o21ai_1 _10400_ (.B1(_04449_),
    .VDD(VPWR),
    .Y(_04450_),
    .VSS(VGND),
    .A1(_04411_),
    .A2(_04448_));
 sg13g2_inv_1 _10401_ (.VDD(VPWR),
    .Y(_04451_),
    .A(_04397_),
    .VSS(VGND));
 sg13g2_nor2_1 _10402_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[8] ),
    .B(_04390_),
    .Y(_04452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10403_ (.A(_04452_),
    .B(_04392_),
    .Y(_04453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10404_ (.VDD(VPWR),
    .Y(_04454_),
    .A(_04453_),
    .VSS(VGND));
 sg13g2_nor2_1 _10405_ (.A(_04451_),
    .B(_04454_),
    .Y(_04455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _10406_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_04455_),
    .C1(_04396_),
    .B1(_04450_),
    .A1(_04392_),
    .Y(_04456_),
    .A2(_04397_));
 sg13g2_nor2_1 _10407_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[10] ),
    .B(_02457_),
    .Y(_04457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10408_ (.VDD(VPWR),
    .Y(_04458_),
    .A(_04457_),
    .VSS(VGND));
 sg13g2_nor2_1 _10409_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_b[10] ),
    .B(_02259_),
    .Y(_04459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _10410_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_04459_),
    .Y(_04460_),
    .A2(_04458_),
    .A1(_04456_));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10412_ (.VDD(VPWR),
    .Y(_04462_),
    .A(\fp16_sum_pipe.reg2en.q[0] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _10413_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04460_),
    .A2(_02177_),
    .Y(_04463_),
    .B1(_04462_));
 sg13g2_o21ai_1 _10414_ (.B1(_04463_),
    .VDD(VPWR),
    .Y(_04464_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.op_sign_logic0.s_a ),
    .A2(_04460_));
 sg13g2_o21ai_1 _10415_ (.B1(_04464_),
    .VDD(VPWR),
    .Y(_01173_),
    .VSS(VGND),
    .A1(net1846),
    .A2(_04389_));
 sg13g2_inv_4 _10416_ (.A(net1838),
    .Y(_04465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10417_ (.Y(_04466_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[10] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10418_ (.B1(\fp16_sum_pipe.reg2en.q[0] ),
    .VDD(VPWR),
    .Y(_04467_),
    .VSS(VGND),
    .A1(_04466_),
    .A2(_04384_));
 sg13g2_nor2_1 _10419_ (.A(_04459_),
    .B(_04457_),
    .Y(_04468_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10420_ (.Y(_04469_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[9] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10421_ (.VDD(VPWR),
    .Y(_04470_),
    .A(_04469_),
    .VSS(VGND));
 sg13g2_nand2_1 _10422_ (.Y(_04471_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[7] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10423_ (.VDD(VPWR),
    .Y(_04472_),
    .A(_04471_),
    .VSS(VGND));
 sg13g2_nand2_1 _10424_ (.Y(_04473_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[0] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10425_ (.Y(_04474_),
    .A(_04412_),
    .B(_04416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _10426_ (.Y(_04475_),
    .B(_04474_),
    .A_N(_04473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10427_ (.Y(_04476_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[1] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10428_ (.Y(_04477_),
    .A(_04475_),
    .B(_04476_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10429_ (.VDD(VPWR),
    .Y(_04478_),
    .A(_04423_),
    .VSS(VGND));
 sg13g2_nand2_1 _10430_ (.Y(_04479_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[2] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10431_ (.VDD(VPWR),
    .Y(_04480_),
    .A(_04479_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10432_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04477_),
    .A2(_04478_),
    .Y(_04481_),
    .B1(_04480_));
 sg13g2_nand2_1 _10433_ (.Y(_04482_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[3] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10434_ (.B1(_04482_),
    .VDD(VPWR),
    .Y(_04483_),
    .VSS(VGND),
    .A1(_04428_),
    .A2(_04481_));
 sg13g2_nand2_1 _10435_ (.Y(_04484_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[4] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10436_ (.VDD(VPWR),
    .Y(_04485_),
    .A(_04484_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04483_),
    .A2(_04437_),
    .Y(_04486_),
    .B1(_04485_));
 sg13g2_nand2_1 _10438_ (.Y(_04487_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[5] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10439_ (.B1(_04487_),
    .VDD(VPWR),
    .Y(_04488_),
    .VSS(VGND),
    .A1(_04442_),
    .A2(_04486_));
 sg13g2_nand2_1 _10440_ (.Y(_04489_),
    .A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[6] ),
    .B(\fp16_sum_pipe.op_sign_logic0.mantisa_b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10441_ (.VDD(VPWR),
    .Y(_04490_),
    .A(_04489_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10442_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04488_),
    .A2(_04409_),
    .Y(_04491_),
    .B1(_04490_));
 sg13g2_nor2_1 _10443_ (.A(_04384_),
    .B(_04491_),
    .Y(_04492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10444_ (.Y(_04493_),
    .B1(_04403_),
    .B2(_04492_),
    .A2(_04472_),
    .A1(net1736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10445_ (.B(\fp16_sum_pipe.op_sign_logic0.mantisa_a[8] ),
    .C(\fp16_sum_pipe.op_sign_logic0.mantisa_b[8] ),
    .A(net1736),
    .Y(_04494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10446_ (.B1(_04494_),
    .VDD(VPWR),
    .Y(_04495_),
    .VSS(VGND),
    .A1(_04453_),
    .A2(_04493_));
 sg13g2_a22oi_1 _10447_ (.Y(_04496_),
    .B1(_04451_),
    .B2(_04495_),
    .A2(_04470_),
    .A1(_04386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10448_ (.A(_04468_),
    .B(_04496_),
    .Y(_04497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10449_ (.A(_04467_),
    .B(_04497_),
    .Y(_04498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10450_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04462_),
    .A2(_04465_),
    .Y(_01172_),
    .B1(_04498_));
 sg13g2_inv_1 _10451_ (.VDD(VPWR),
    .Y(_04499_),
    .A(_04468_),
    .VSS(VGND));
 sg13g2_nor2_1 _10452_ (.A(\fp16_sum_pipe.op_sign_logic0.mantisa_a[0] ),
    .B(_04413_),
    .Y(_04500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _10453_ (.Y(_04501_),
    .B(_04414_),
    .A_N(_04500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10454_ (.A(_04474_),
    .B(_04501_),
    .C(_04429_),
    .Y(_04502_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10455_ (.A(_04499_),
    .B(_04451_),
    .C(_04454_),
    .Y(_04503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _10456_ (.B(_04503_),
    .C(_04410_),
    .A(_04502_),
    .Y(_04504_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04444_));
 sg13g2_nand2_1 _10457_ (.Y(_04505_),
    .A(_04504_),
    .B(_04458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10458_ (.B1(_04412_),
    .VDD(VPWR),
    .Y(_04506_),
    .VSS(VGND),
    .A1(_04500_),
    .A2(_04417_));
 sg13g2_a21oi_1 _10459_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04506_),
    .A2(_04423_),
    .Y(_04507_),
    .B1(_04422_));
 sg13g2_inv_1 _10460_ (.VDD(VPWR),
    .Y(_04508_),
    .A(_04507_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10461_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04508_),
    .A2(_04426_),
    .Y(_04509_),
    .B1(_04425_));
 sg13g2_inv_1 _10462_ (.VDD(VPWR),
    .Y(_04510_),
    .A(_04509_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10463_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04510_),
    .A2(_04436_),
    .Y(_04511_),
    .B1(_04435_));
 sg13g2_inv_1 _10464_ (.VDD(VPWR),
    .Y(_04512_),
    .A(_04511_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10465_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04512_),
    .A2(_04440_),
    .Y(_04513_),
    .B1(_04439_));
 sg13g2_a21oi_1 _10466_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04405_),
    .A2(_04400_),
    .Y(_04514_),
    .B1(_04399_));
 sg13g2_o21ai_1 _10467_ (.B1(_04514_),
    .VDD(VPWR),
    .Y(_04515_),
    .VSS(VGND),
    .A1(_04411_),
    .A2(_04513_));
 sg13g2_a221oi_1 _10468_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_04455_),
    .C1(_04394_),
    .B1(_04515_),
    .A1(_04452_),
    .Y(_04516_),
    .A2(_04397_));
 sg13g2_nor2_1 _10469_ (.A(_04505_),
    .B(_04516_),
    .Y(_04517_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10470_ (.B1(_04384_),
    .VDD(VPWR),
    .Y(_04518_),
    .VSS(VGND),
    .A1(_04459_),
    .A2(_04456_));
 sg13g2_o21ai_1 _10471_ (.B1(_04496_),
    .VDD(VPWR),
    .Y(_04519_),
    .VSS(VGND),
    .A1(_04517_),
    .A2(_04518_));
 sg13g2_xnor2_1 _10472_ (.Y(_04520_),
    .A(_04499_),
    .B(_04519_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10473_ (.A(net1847),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[10] ),
    .Y(_04521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10474_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04520_),
    .A2(net1847),
    .Y(_01171_),
    .B1(_04521_));
 sg13g2_inv_1 _10475_ (.VDD(VPWR),
    .Y(_04522_),
    .A(_04450_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10476_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04522_),
    .A2(_04391_),
    .Y(_04523_),
    .B1(_04452_));
 sg13g2_a21oi_1 _10477_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04515_),
    .A2(_04453_),
    .Y(_04524_),
    .B1(_04452_));
 sg13g2_nor2_1 _10478_ (.A(_04460_),
    .B(_04524_),
    .Y(_04525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10479_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1673),
    .A2(_04523_),
    .Y(_04526_),
    .B1(_04525_));
 sg13g2_a21oi_1 _10480_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04384_),
    .A2(_04526_),
    .Y(_04527_),
    .B1(_04495_));
 sg13g2_xnor2_1 _10481_ (.Y(_04528_),
    .A(_04397_),
    .B(_04527_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10482_ (.A(net1847),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[9] ),
    .Y(_04529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10483_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04528_),
    .A2(net1847),
    .Y(_01170_),
    .B1(_04529_));
 sg13g2_inv_1 _10484_ (.VDD(VPWR),
    .Y(_04530_),
    .A(_04460_),
    .VSS(VGND));
 sg13g2_nor2_1 _10485_ (.A(_04522_),
    .B(_04530_),
    .Y(_04531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _10486_ (.A2(_04515_),
    .A1(net1670),
    .B1(net1736),
    .X(_04532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10487_ (.B1(_04493_),
    .VDD(VPWR),
    .Y(_04533_),
    .VSS(VGND),
    .A1(_04531_),
    .A2(_04532_));
 sg13g2_xnor2_1 _10488_ (.Y(_04534_),
    .A(_04454_),
    .B(_04533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10489_ (.A(net1847),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[8] ),
    .Y(_04535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10490_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04534_),
    .A2(net1847),
    .Y(_01169_),
    .B1(_04535_));
 sg13g2_a21oi_1 _10491_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04447_),
    .A2(_04408_),
    .Y(_04536_),
    .B1(_04407_));
 sg13g2_nor2_1 _10492_ (.A(_04536_),
    .B(net1670),
    .Y(_04537_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10493_ (.VDD(VPWR),
    .Y(_04538_),
    .A(_04513_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10494_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04538_),
    .A2(_04408_),
    .Y(_04539_),
    .B1(_04405_));
 sg13g2_o21ai_1 _10495_ (.B1(_04384_),
    .VDD(VPWR),
    .Y(_04540_),
    .VSS(VGND),
    .A1(_04539_),
    .A2(net1673));
 sg13g2_inv_1 _10496_ (.VDD(VPWR),
    .Y(_04541_),
    .A(_04492_),
    .VSS(VGND));
 sg13g2_o21ai_1 _10497_ (.B1(_04541_),
    .VDD(VPWR),
    .Y(_04542_),
    .VSS(VGND),
    .A1(_04537_),
    .A2(_04540_));
 sg13g2_xnor2_1 _10498_ (.Y(_04543_),
    .A(_04403_),
    .B(_04542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10499_ (.A(net1847),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[7] ),
    .Y(_04544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10500_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04543_),
    .A2(net1848),
    .Y(_01168_),
    .B1(_04544_));
 sg13g2_nand2_1 _10501_ (.Y(_04545_),
    .A(net1670),
    .B(_04538_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10502_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1673),
    .A2(_04447_),
    .Y(_04546_),
    .B1(net1736));
 sg13g2_a22oi_1 _10503_ (.Y(_04547_),
    .B1(_04545_),
    .B2(_04546_),
    .A2(_04488_),
    .A1(net1736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10504_ (.Y(_04548_),
    .A(_04408_),
    .B(_04547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10505_ (.A(net1848),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[6] ),
    .Y(_04549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10506_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04548_),
    .A2(net1848),
    .Y(_01167_),
    .B1(_04549_));
 sg13g2_nand2_1 _10507_ (.Y(_04550_),
    .A(net1670),
    .B(_04512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04431_),
    .A2(_04436_),
    .Y(_04551_),
    .B1(_04433_));
 sg13g2_nand2b_1 _10509_ (.Y(_04552_),
    .B(net1673),
    .A_N(_04551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10510_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04550_),
    .A2(_04552_),
    .Y(_04553_),
    .B1(net1736));
 sg13g2_a21oi_1 _10511_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1736),
    .A2(_04486_),
    .Y(_04554_),
    .B1(_04553_));
 sg13g2_xnor2_1 _10512_ (.Y(_04555_),
    .A(_04443_),
    .B(_04554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10513_ (.A(net1848),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[5] ),
    .Y(_04556_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10514_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04555_),
    .A2(net1848),
    .Y(_01166_),
    .B1(_04556_));
 sg13g2_nand2_1 _10515_ (.Y(_04557_),
    .A(net1673),
    .B(_04431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10516_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1670),
    .A2(_04510_),
    .Y(_04558_),
    .B1(net1737));
 sg13g2_a22oi_1 _10517_ (.Y(_04559_),
    .B1(_04557_),
    .B2(_04558_),
    .A2(_04483_),
    .A1(net1737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10518_ (.Y(_04560_),
    .A(_04436_),
    .B(_04559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10519_ (.A(net1848),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .Y(_04561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10520_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04560_),
    .A2(net1848),
    .Y(_01165_),
    .B1(_04561_));
 sg13g2_inv_1 _10521_ (.VDD(VPWR),
    .Y(_04562_),
    .A(_04481_),
    .VSS(VGND));
 sg13g2_nor2_1 _10522_ (.A(_04478_),
    .B(_04418_),
    .Y(_04563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10523_ (.B1(net1673),
    .VDD(VPWR),
    .Y(_04564_),
    .VSS(VGND),
    .A1(_04420_),
    .A2(_04563_));
 sg13g2_a21oi_1 _10524_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1670),
    .A2(_04508_),
    .Y(_04565_),
    .B1(net1737));
 sg13g2_a22oi_1 _10525_ (.Y(_04566_),
    .B1(_04564_),
    .B2(_04565_),
    .A2(_04562_),
    .A1(net1737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10526_ (.Y(_04567_),
    .A(_04428_),
    .B(_04566_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10527_ (.A(net1849),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .Y(_04568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10528_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04567_),
    .A2(net1849),
    .Y(_01164_),
    .B1(_04568_));
 sg13g2_nand2b_1 _10529_ (.Y(_04569_),
    .B(net1673),
    .A_N(_04418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10530_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1670),
    .A2(_04506_),
    .Y(_04570_),
    .B1(net1737));
 sg13g2_a22oi_1 _10531_ (.Y(_04571_),
    .B1(_04569_),
    .B2(_04570_),
    .A2(_04477_),
    .A1(net1737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10532_ (.Y(_04572_),
    .A(_04423_),
    .B(_04571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10533_ (.A(net1849),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[2] ),
    .Y(_04573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10534_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04572_),
    .A2(net1849),
    .Y(_01163_),
    .B1(_04573_));
 sg13g2_nand2b_1 _10535_ (.Y(_04574_),
    .B(net1673),
    .A_N(_04414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10536_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1670),
    .A2(_04500_),
    .Y(_04575_),
    .B1(net1737));
 sg13g2_a22oi_1 _10537_ (.Y(_04576_),
    .B1(_04574_),
    .B2(_04575_),
    .A2(_04473_),
    .A1(net1737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10538_ (.Y(_04577_),
    .A(_04474_),
    .B(_04576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10539_ (.A(net1849),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[1] ),
    .Y(_04578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10540_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04577_),
    .A2(net1849),
    .Y(_01162_),
    .B1(_04578_));
 sg13g2_inv_1 _10541_ (.VDD(VPWR),
    .Y(_04579_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10542_ (.Y(_04580_),
    .A(_04501_),
    .B(net1849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10543_ (.B1(_04580_),
    .VDD(VPWR),
    .Y(_01161_),
    .VSS(VGND),
    .A1(net1849),
    .A2(_04579_));
 sg13g2_inv_2 _10544_ (.Y(_04581_),
    .A(\fp16_sum_pipe.add_renorm0.exp[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10545_ (.Y(_04582_),
    .A(\fp16_sum_pipe.seg_reg0.q[29] ),
    .B(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10546_ (.B1(_04582_),
    .VDD(VPWR),
    .Y(_01160_),
    .VSS(VGND),
    .A1(net1846),
    .A2(_04581_));
 sg13g2_inv_1 _10547_ (.VDD(VPWR),
    .Y(_04583_),
    .A(\fp16_sum_pipe.add_renorm0.exp[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10548_ (.Y(_04584_),
    .A(\fp16_sum_pipe.seg_reg0.q[28] ),
    .B(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10549_ (.B1(_04584_),
    .VDD(VPWR),
    .Y(_01159_),
    .VSS(VGND),
    .A1(net1846),
    .A2(_04583_));
 sg13g2_inv_2 _10550_ (.Y(_04585_),
    .A(\fp16_sum_pipe.add_renorm0.exp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10551_ (.Y(_04586_),
    .A(\fp16_sum_pipe.seg_reg0.q[27] ),
    .B(net1846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10552_ (.B1(_04586_),
    .VDD(VPWR),
    .Y(_01158_),
    .VSS(VGND),
    .A1(net1846),
    .A2(_04585_));
 sg13g2_inv_2 _10553_ (.Y(_04587_),
    .A(\fp16_sum_pipe.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10554_ (.Y(_04588_),
    .A(\fp16_sum_pipe.seg_reg0.q[26] ),
    .B(net1846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10555_ (.B1(_04588_),
    .VDD(VPWR),
    .Y(_01157_),
    .VSS(VGND),
    .A1(net1846),
    .A2(_04587_));
 sg13g2_inv_2 _10556_ (.Y(_04589_),
    .A(\fp16_sum_pipe.add_renorm0.exp[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10557_ (.Y(_04590_),
    .A(\fp16_sum_pipe.seg_reg0.q[25] ),
    .B(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10558_ (.B1(_04590_),
    .VDD(VPWR),
    .Y(_01156_),
    .VSS(VGND),
    .A1(net1845),
    .A2(_04589_));
 sg13g2_inv_1 _10559_ (.VDD(VPWR),
    .Y(_04591_),
    .A(\fp16_sum_pipe.add_renorm0.exp[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10560_ (.Y(_04592_),
    .A(\fp16_sum_pipe.seg_reg0.q[24] ),
    .B(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10561_ (.B1(_04592_),
    .VDD(VPWR),
    .Y(_01155_),
    .VSS(VGND),
    .A1(net1844),
    .A2(_04591_));
 sg13g2_inv_1 _10562_ (.VDD(VPWR),
    .Y(_04593_),
    .A(\fp16_sum_pipe.add_renorm0.exp[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10563_ (.Y(_04594_),
    .A(\fp16_sum_pipe.seg_reg0.q[23] ),
    .B(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10564_ (.B1(_04594_),
    .VDD(VPWR),
    .Y(_01154_),
    .VSS(VGND),
    .A1(net1844),
    .A2(_04593_));
 sg13g2_inv_1 _10565_ (.VDD(VPWR),
    .Y(_04595_),
    .A(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10566_ (.Y(_04596_),
    .A(\fp16_sum_pipe.seg_reg0.q[22] ),
    .B(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10567_ (.B1(_04596_),
    .VDD(VPWR),
    .Y(_01153_),
    .VSS(VGND),
    .A1(net1844),
    .A2(_04595_));
 sg13g2_nor2_1 _10568_ (.A(\fp16_sum_pipe.exp_mant_logic0.a[15] ),
    .B(net1931),
    .Y(_04597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10569_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03327_),
    .A2(net1931),
    .Y(_01152_),
    .B1(_04597_));
 sg13g2_nand2_1 _10570_ (.Y(_04598_),
    .A(\acc_sub.x2[14] ),
    .B(net1925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10571_ (.B1(_04598_),
    .VDD(VPWR),
    .Y(_01151_),
    .VSS(VGND),
    .A1(net1925),
    .A2(_02238_));
 sg13g2_nand2_1 _10572_ (.Y(_04599_),
    .A(\acc_sub.x2[13] ),
    .B(net1931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10573_ (.B1(_04599_),
    .VDD(VPWR),
    .Y(_01150_),
    .VSS(VGND),
    .A1(net1931),
    .A2(_02186_));
 sg13g2_nand2_1 _10574_ (.Y(_04600_),
    .A(\acc_sub.x2[12] ),
    .B(net1924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10575_ (.B1(_04600_),
    .VDD(VPWR),
    .Y(_01149_),
    .VSS(VGND),
    .A1(net1926),
    .A2(_02197_));
 sg13g2_nand2_1 _10576_ (.Y(_04601_),
    .A(\acc_sub.x2[11] ),
    .B(net1924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10577_ (.B1(_04601_),
    .VDD(VPWR),
    .Y(_01148_),
    .VSS(VGND),
    .A1(net1926),
    .A2(_02192_));
 sg13g2_nand2_1 _10578_ (.Y(_04602_),
    .A(\acc_sub.x2[10] ),
    .B(net1931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10579_ (.B1(_04602_),
    .VDD(VPWR),
    .Y(_01147_),
    .VSS(VGND),
    .A1(net1930),
    .A2(_02203_));
 sg13g2_nand2_1 _10580_ (.Y(_04603_),
    .A(\acc_sub.x2[9] ),
    .B(net1925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10581_ (.B1(_04603_),
    .VDD(VPWR),
    .Y(_01146_),
    .VSS(VGND),
    .A1(net1930),
    .A2(_02208_));
 sg13g2_nand2_1 _10582_ (.Y(_04604_),
    .A(\acc_sub.x2[8] ),
    .B(net1926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10583_ (.B1(_04604_),
    .VDD(VPWR),
    .Y(_01145_),
    .VSS(VGND),
    .A1(net1932),
    .A2(_02264_));
 sg13g2_nand2_1 _10584_ (.Y(_04605_),
    .A(\acc_sub.x2[7] ),
    .B(net1931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10585_ (.B1(_04605_),
    .VDD(VPWR),
    .Y(_01144_),
    .VSS(VGND),
    .A1(net1932),
    .A2(_02218_));
 sg13g2_nand2_1 _10586_ (.Y(_04606_),
    .A(\acc_sub.x2[6] ),
    .B(net1932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10587_ (.B1(_04606_),
    .VDD(VPWR),
    .Y(_01143_),
    .VSS(VGND),
    .A1(net1927),
    .A2(_02267_));
 sg13g2_nand2_1 _10588_ (.Y(_04607_),
    .A(\acc_sub.x2[5] ),
    .B(net1934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10589_ (.B1(_04607_),
    .VDD(VPWR),
    .Y(_01142_),
    .VSS(VGND),
    .A1(net1934),
    .A2(_02260_));
 sg13g2_nand2_1 _10590_ (.Y(_04608_),
    .A(\acc_sub.x2[4] ),
    .B(net1927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10591_ (.B1(_04608_),
    .VDD(VPWR),
    .Y(_01141_),
    .VSS(VGND),
    .A1(net1927),
    .A2(_02261_));
 sg13g2_nand2_1 _10592_ (.Y(_04609_),
    .A(\acc_sub.x2[3] ),
    .B(net1934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10593_ (.B1(_04609_),
    .VDD(VPWR),
    .Y(_01140_),
    .VSS(VGND),
    .A1(net1934),
    .A2(_02268_));
 sg13g2_nand2_1 _10594_ (.Y(_04610_),
    .A(\acc_sub.x2[2] ),
    .B(net1934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10595_ (.B1(_04610_),
    .VDD(VPWR),
    .Y(_01139_),
    .VSS(VGND),
    .A1(net1933),
    .A2(_02269_));
 sg13g2_nand2_1 _10596_ (.Y(_04611_),
    .A(\acc_sub.x2[1] ),
    .B(net1933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10597_ (.B1(_04611_),
    .VDD(VPWR),
    .Y(_01138_),
    .VSS(VGND),
    .A1(net1934),
    .A2(_02262_));
 sg13g2_nand2_1 _10598_ (.Y(_04612_),
    .A(\acc_sub.x2[0] ),
    .B(net1933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10599_ (.B1(_04612_),
    .VDD(VPWR),
    .Y(_01137_),
    .VSS(VGND),
    .A1(net1934),
    .A2(_02270_));
 sg13g2_inv_1 _10600_ (.VDD(VPWR),
    .Y(_04613_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10601_ (.Y(_04614_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .B(\fp16_res_pipe.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10602_ (.B1(_04614_),
    .VDD(VPWR),
    .Y(_04615_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .A2(_04613_));
 sg13g2_inv_1 _10603_ (.VDD(VPWR),
    .Y(_04616_),
    .A(net1823),
    .VSS(VGND));
 sg13g2_nand2_1 _10604_ (.Y(_04617_),
    .A(net1823),
    .B(\fp16_res_pipe.add_renorm0.mantisa[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10605_ (.VDD(VPWR),
    .Y(_04618_),
    .A(_04617_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10606_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04616_),
    .A2(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .Y(_04619_),
    .B1(_04618_));
 sg13g2_inv_1 _10607_ (.VDD(VPWR),
    .Y(_04620_),
    .A(_04619_),
    .VSS(VGND));
 sg13g2_inv_2 _10608_ (.Y(_04621_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10609_ (.Y(_04622_),
    .A(_04621_),
    .B(net1826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10610_ (.B1(_04622_),
    .VDD(VPWR),
    .Y(_04623_),
    .VSS(VGND),
    .A1(net1826),
    .A2(\fp16_res_pipe.add_renorm0.mantisa[4] ));
 sg13g2_inv_1 _10611_ (.VDD(VPWR),
    .Y(_04624_),
    .A(_04623_),
    .VSS(VGND));
 sg13g2_nand2_1 _10612_ (.Y(_04625_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .B(\fp16_res_pipe.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10613_ (.B1(_04625_),
    .VDD(VPWR),
    .Y(_04626_),
    .VSS(VGND),
    .A1(net1826),
    .A2(_04621_));
 sg13g2_nand3_1 _10614_ (.B(_04624_),
    .C(_04626_),
    .A(_04620_),
    .Y(_04627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10615_ (.VDD(VPWR),
    .Y(_04628_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10616_ (.A(net1823),
    .B(\fp16_res_pipe.add_renorm0.mantisa[2] ),
    .Y(_04629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10617_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1823),
    .A2(_04628_),
    .Y(_04630_),
    .B1(_04629_));
 sg13g2_inv_1 _10618_ (.VDD(VPWR),
    .Y(_04631_),
    .A(_04630_),
    .VSS(VGND));
 sg13g2_nor2_1 _10619_ (.A(_04619_),
    .B(_04631_),
    .Y(_04632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10620_ (.VDD(VPWR),
    .Y(_04633_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[2] ),
    .VSS(VGND));
 sg13g2_a22oi_1 _10621_ (.Y(_04634_),
    .B1(_04616_),
    .B2(_03572_),
    .A2(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .A1(_04633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10622_ (.A(\fp16_res_pipe.add_renorm0.mantisa[1] ),
    .B(_04629_),
    .C(_04634_),
    .Y(_04635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10623_ (.A(_04631_),
    .B(_04635_),
    .Y(_04636_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10624_ (.A(_04632_),
    .B(_04636_),
    .Y(_04637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10625_ (.A(_04627_),
    .B(_04637_),
    .Y(_04638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10626_ (.Y(_04639_),
    .A(_04615_),
    .B(_04638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10627_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03565_),
    .A2(_03572_),
    .Y(_04640_),
    .B1(_04633_));
 sg13g2_nand2_1 _10628_ (.Y(_04641_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .B(\fp16_res_pipe.add_renorm0.mantisa[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10629_ (.B1(_04641_),
    .VDD(VPWR),
    .Y(_04642_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .A2(_04640_));
 sg13g2_buf_2 place1744 (.A(_01496_),
    .X(net1744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10631_ (.VDD(VPWR),
    .Y(_04644_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[7] ),
    .VSS(VGND));
 sg13g2_nand4_1 _10632_ (.B(\fp16_res_pipe.add_renorm0.mantisa[4] ),
    .C(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .A(\fp16_res_pipe.add_renorm0.mantisa[5] ),
    .Y(_04645_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\fp16_res_pipe.add_renorm0.mantisa[2] ));
 sg13g2_nor2_1 _10633_ (.A(_04613_),
    .B(_04645_),
    .Y(_04646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10634_ (.Y(_04647_),
    .A(_04644_),
    .B(_04646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1752 (.A(net1751),
    .X(net1752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10636_ (.VDD(VPWR),
    .Y(_04649_),
    .A(_04647_),
    .VSS(VGND));
 sg13g2_nand3_1 _10637_ (.B(\fp16_res_pipe.add_renorm0.mantisa[8] ),
    .C(\fp16_res_pipe.add_renorm0.mantisa[7] ),
    .A(_04646_),
    .Y(_04650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10638_ (.VDD(VPWR),
    .Y(_04651_),
    .A(_04650_),
    .VSS(VGND));
 sg13g2_nand2_2 _10639_ (.Y(_04652_),
    .A(_04651_),
    .B(\fp16_res_pipe.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10640_ (.VDD(VPWR),
    .Y(_04653_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[10] ),
    .VSS(VGND));
 sg13g2_nand2_2 _10641_ (.Y(_04654_),
    .A(_04652_),
    .B(_04653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10642_ (.VDD(VPWR),
    .Y(_04655_),
    .A(_04652_),
    .VSS(VGND));
 sg13g2_inv_1 _10643_ (.VDD(VPWR),
    .Y(_04656_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _10644_ (.Y(_04657_),
    .A(_04650_),
    .B(_04656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _10645_ (.A(_04655_),
    .B_N(_04657_),
    .Y(_04658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1713 (.A(_06907_),
    .X(net1713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10647_ (.A(_04654_),
    .B(_04658_),
    .Y(_04660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _10648_ (.A2(\fp16_res_pipe.add_renorm0.mantisa[7] ),
    .A1(_04646_),
    .B1(\fp16_res_pipe.add_renorm0.mantisa[8] ),
    .X(_04661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10649_ (.A(_04661_),
    .B(_04650_),
    .X(_04662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout95 (.A(net96),
    .X(net95),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10651_ (.Y(_04664_),
    .A(_04662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10652_ (.Y(_04665_),
    .A(_04660_),
    .B(_04664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10653_ (.A(_04649_),
    .B(_04665_),
    .Y(_04666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10654_ (.VDD(VPWR),
    .Y(_04667_),
    .A(_04666_),
    .VSS(VGND));
 sg13g2_nor2_1 _10655_ (.A(_04642_),
    .B(_04667_),
    .Y(_04668_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1750 (.A(net1749),
    .X(net1750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _10657_ (.A(_04654_),
    .B(_04658_),
    .C(_04664_),
    .Y(_04670_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1692 (.A(_02244_),
    .X(net1692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10659_ (.Y(_04672_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[4] ),
    .B(_04641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1753 (.A(net1752),
    .X(net1753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10661_ (.Y(_04674_),
    .A(_04670_),
    .B(_04672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10662_ (.Y(_04675_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[6] ),
    .B(_04645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout69 (.A(net70),
    .X(net69),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10664_ (.Y(_04677_),
    .A(net1710),
    .B(_04675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10665_ (.VDD(VPWR),
    .Y(_04678_),
    .A(_04658_),
    .VSS(VGND));
 sg13g2_nor2_2 _10666_ (.A(_04654_),
    .B(_04678_),
    .Y(_04679_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _10667_ (.A(_04641_),
    .B_N(\fp16_res_pipe.add_renorm0.mantisa[4] ),
    .Y(_04680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10668_ (.Y(_04681_),
    .A(_04621_),
    .B(_04680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout85 (.A(net86),
    .X(net85),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10670_ (.Y(_04683_),
    .A(_04679_),
    .B(_04681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10671_ (.B(_04677_),
    .C(_04683_),
    .A(_04674_),
    .Y(_04684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10672_ (.B1(net1822),
    .VDD(VPWR),
    .Y(_04685_),
    .VSS(VGND),
    .A1(_04668_),
    .A2(_04684_));
 sg13g2_o21ai_1 _10673_ (.B1(_04685_),
    .VDD(VPWR),
    .Y(_04686_),
    .VSS(VGND),
    .A1(net1822),
    .A2(_04639_));
 sg13g2_nand2_1 _10674_ (.Y(_04687_),
    .A(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .B(\fp16_res_pipe.add_renorm0.mantisa[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10675_ (.B1(_04687_),
    .VDD(VPWR),
    .Y(_04688_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .A2(_04644_));
 sg13g2_inv_1 _10676_ (.VDD(VPWR),
    .Y(_04689_),
    .A(_04688_),
    .VSS(VGND));
 sg13g2_nand2_1 _10677_ (.Y(_04690_),
    .A(_04638_),
    .B(_04615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10678_ (.Y(_04691_),
    .A(_04689_),
    .B(_04690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10679_ (.A(_04647_),
    .B(_04658_),
    .Y(_04692_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10680_ (.B(_04664_),
    .C(_04675_),
    .A(_04692_),
    .Y(_04693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10681_ (.A(net1710),
    .B(_04693_),
    .Y(_04694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10682_ (.Y(_04695_),
    .A(_04642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10683_ (.Y(_04696_),
    .A(_04694_),
    .B(_04695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10684_ (.Y(_04697_),
    .B1(_04675_),
    .B2(_04679_),
    .A2(net1710),
    .A1(_04647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10685_ (.Y(_04698_),
    .A(_04666_),
    .B(_04672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10686_ (.Y(_04699_),
    .A(_04670_),
    .B(_04681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _10687_ (.B(_04697_),
    .C(_04698_),
    .A(_04696_),
    .Y(_04700_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04699_));
 sg13g2_nand2_1 _10688_ (.Y(_04701_),
    .A(_04700_),
    .B(net1822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10689_ (.B1(_04701_),
    .VDD(VPWR),
    .Y(_04702_),
    .VSS(VGND),
    .A1(net1822),
    .A2(_04691_));
 sg13g2_a22oi_1 _10690_ (.Y(_04703_),
    .B1(_04695_),
    .B2(_04679_),
    .A2(_04672_),
    .A1(net1710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10691_ (.VDD(VPWR),
    .Y(_04704_),
    .A(_04632_),
    .VSS(VGND));
 sg13g2_nor2_1 _10692_ (.A(_04623_),
    .B(_04704_),
    .Y(_04705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10693_ (.Y(_04706_),
    .A(_04704_),
    .B(_04623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _10694_ (.B(_03359_),
    .C(_04706_),
    .Y(_04707_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_04705_));
 sg13g2_o21ai_1 _10695_ (.B1(_04707_),
    .VDD(VPWR),
    .Y(_04708_),
    .VSS(VGND),
    .A1(net1771),
    .A2(_04703_));
 sg13g2_nand2_1 _10696_ (.Y(_04709_),
    .A(net1826),
    .B(\fp16_res_pipe.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10697_ (.B1(_04709_),
    .VDD(VPWR),
    .Y(_04710_),
    .VSS(VGND),
    .A1(net1826),
    .A2(_03512_));
 sg13g2_and3_1 _10698_ (.X(_04711_),
    .A(_04710_),
    .B(_04688_),
    .C(_04615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10699_ (.Y(_04712_),
    .A(_04638_),
    .B(_04711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10700_ (.Y(_04713_),
    .A(net1826),
    .B(\fp16_res_pipe.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10701_ (.B1(_04713_),
    .VDD(VPWR),
    .Y(_04714_),
    .VSS(VGND),
    .A1(net1826),
    .A2(_04656_));
 sg13g2_inv_1 _10702_ (.VDD(VPWR),
    .Y(_04715_),
    .A(_04714_),
    .VSS(VGND));
 sg13g2_nand3b_1 _10703_ (.B(_04711_),
    .C(_04714_),
    .Y(_04716_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_04627_));
 sg13g2_nor2_1 _10704_ (.A(_04637_),
    .B(_04716_),
    .Y(_04717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _10705_ (.A2(_04715_),
    .A1(_04712_),
    .B1(_04717_),
    .X(_04718_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _10706_ (.Y(_04719_),
    .B(_04681_),
    .A_N(_04675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _10707_ (.A(_04647_),
    .B(_04719_),
    .C(_04665_),
    .Y(_04720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10708_ (.Y(_04721_),
    .B1(_04672_),
    .B2(_04720_),
    .A2(_04681_),
    .A1(_04694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10709_ (.A(_04647_),
    .B(_04665_),
    .Y(_04722_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10710_ (.A(_04681_),
    .B(_04675_),
    .Y(_04723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10711_ (.B(_04672_),
    .C(_04723_),
    .A(_04722_),
    .Y(_04724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1694 (.A(net1693),
    .X(net1694),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10713_ (.VDD(VPWR),
    .Y(_04726_),
    .A(_04724_),
    .VSS(VGND));
 sg13g2_nand2_1 _10714_ (.Y(_04727_),
    .A(_04726_),
    .B(_04695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10715_ (.B1(_04658_),
    .VDD(VPWR),
    .Y(_04728_),
    .VSS(VGND),
    .A1(net1710),
    .A2(_04662_));
 sg13g2_a22oi_1 _10716_ (.Y(_04729_),
    .B1(_04675_),
    .B2(_04666_),
    .A2(_04670_),
    .A1(_04647_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _10717_ (.B(_04727_),
    .C(_04728_),
    .A(_04721_),
    .Y(_04730_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04729_));
 sg13g2_nand2_1 _10718_ (.Y(_04731_),
    .A(_04730_),
    .B(net1822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10719_ (.B1(_04731_),
    .VDD(VPWR),
    .Y(_04732_),
    .VSS(VGND),
    .A1(net1821),
    .A2(_04718_));
 sg13g2_nor4_1 _10720_ (.A(_04686_),
    .B(_04702_),
    .C(_04708_),
    .D(_04732_),
    .Y(_04733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _10721_ (.A(_04681_),
    .B(_04672_),
    .C(_04642_),
    .D(_04675_),
    .Y(_04734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _10722_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_04720_),
    .Y(_04735_),
    .A2(_04734_),
    .A1(_04722_));
 sg13g2_inv_1 _10723_ (.VDD(VPWR),
    .Y(_04736_),
    .A(_04679_),
    .VSS(VGND));
 sg13g2_nand3_1 _10724_ (.B(_04667_),
    .C(_04736_),
    .A(_04735_),
    .Y(_04737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1674 (.A(_03453_),
    .X(net1674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10726_ (.VDD(VPWR),
    .Y(_04739_),
    .A(_04737_),
    .VSS(VGND));
 sg13g2_inv_2 _10727_ (.Y(_04740_),
    .A(net1710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10728_ (.Y(_04741_),
    .A(_04693_),
    .B(_04740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10729_ (.A(_04670_),
    .B(_04726_),
    .Y(_04742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10730_ (.Y(_04743_),
    .A(_04742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10731_ (.A(_04741_),
    .B(_04743_),
    .Y(_04744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10732_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04739_),
    .A2(_04744_),
    .Y(_04745_),
    .B1(net1771));
 sg13g2_nor2_2 _10733_ (.A(net1824),
    .B(\fp16_res_pipe.add_renorm0.mantisa[10] ),
    .Y(_04746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10734_ (.VDD(VPWR),
    .Y(_04747_),
    .A(_04717_),
    .VSS(VGND));
 sg13g2_nor2_2 _10735_ (.A(_04746_),
    .B(_04747_),
    .Y(_04748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10736_ (.A(_04746_),
    .B(_04630_),
    .Y(_04749_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _10737_ (.B(_04716_),
    .A(_04746_),
    .X(_04750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10738_ (.A(_04750_),
    .B(_04635_),
    .X(_04751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10739_ (.A(_04750_),
    .B(_04636_),
    .X(_04752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _10740_ (.A(_04748_),
    .B(_04749_),
    .C(_04751_),
    .D(_04752_),
    .Y(_04753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10741_ (.B1(net1822),
    .VDD(VPWR),
    .Y(_04754_),
    .VSS(VGND),
    .A1(_04642_),
    .A2(_04740_));
 sg13g2_nor2b_1 _10742_ (.A(_04753_),
    .B_N(_04754_),
    .Y(_04755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10743_ (.Y(_04756_),
    .A(_04626_),
    .B(_04705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10744_ (.B1(_04704_),
    .VDD(VPWR),
    .Y(_04757_),
    .VSS(VGND),
    .A1(_04620_),
    .A2(_04636_));
 sg13g2_nand2_1 _10745_ (.Y(_04758_),
    .A(_04757_),
    .B(net1771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10746_ (.Y(_04759_),
    .A(_04754_),
    .B(_04758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10747_ (.B1(_04759_),
    .VDD(VPWR),
    .Y(_04760_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.seg_reg1.q[21] ),
    .A2(_04756_));
 sg13g2_nor2_1 _10748_ (.A(_04689_),
    .B(_04690_),
    .Y(_04761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10749_ (.B1(_04712_),
    .VDD(VPWR),
    .Y(_04762_),
    .VSS(VGND),
    .A1(_04710_),
    .A2(_04761_));
 sg13g2_a22oi_1 _10750_ (.Y(_04763_),
    .B1(_04695_),
    .B2(_04720_),
    .A2(_04672_),
    .A1(_04694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10751_ (.Y(_04764_),
    .B1(_04647_),
    .B2(_04679_),
    .A2(_04662_),
    .A1(net1710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _10752_ (.Y(_04765_),
    .B1(_04681_),
    .B2(_04666_),
    .A2(_04670_),
    .A1(_04675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10753_ (.B(_04764_),
    .C(_04765_),
    .A(_04763_),
    .Y(_04766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10754_ (.Y(_04767_),
    .A(_04766_),
    .B(net1822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10755_ (.B1(_04767_),
    .VDD(VPWR),
    .Y(_04768_),
    .VSS(VGND),
    .A1(net1822),
    .A2(_04762_));
 sg13g2_nor4_1 _10756_ (.A(_04745_),
    .B(_04755_),
    .C(_04760_),
    .D(_04768_),
    .Y(_04769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10757_ (.Y(_04770_),
    .A(_04733_),
    .B(_04769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10758_ (.Y(_04771_),
    .A(_04770_),
    .B(\fp16_res_pipe.reg3en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _10759_ (.A(net1835),
    .Y(_04772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10760_ (.Y(_04773_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10761_ (.B1(_04773_),
    .VDD(VPWR),
    .Y(_01136_),
    .VSS(VGND),
    .A1(_03367_),
    .A2(_04771_));
 sg13g2_inv_2 _10762_ (.Y(_04774_),
    .A(_04741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10763_ (.A(_04653_),
    .B(_04652_),
    .Y(_04775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout117 (.A(net119),
    .X(net117),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10765_ (.B(\fp16_res_pipe.add_renorm0.exp[1] ),
    .C(\fp16_res_pipe.add_renorm0.exp[0] ),
    .A(\fp16_res_pipe.add_renorm0.exp[2] ),
    .Y(_04777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10766_ (.A(_03582_),
    .B(_04777_),
    .Y(_04778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10767_ (.Y(_04779_),
    .A(_04778_),
    .B(\fp16_res_pipe.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10768_ (.A(_03578_),
    .B(_04779_),
    .Y(_04780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10769_ (.Y(_04781_),
    .A(_04780_),
    .B(\fp16_res_pipe.add_renorm0.exp[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10770_ (.Y(_04782_),
    .A(_03574_),
    .B(_04781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10771_ (.A(\fp16_res_pipe.add_renorm0.exp[7] ),
    .B(net1709),
    .Y(_04783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10772_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1709),
    .A2(_04782_),
    .Y(_04784_),
    .B1(_04783_));
 sg13g2_inv_2 _10773_ (.Y(_04785_),
    .A(_04784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10774_ (.B(\fp16_res_pipe.add_renorm0.mantisa[10] ),
    .C(\fp16_res_pipe.add_renorm0.mantisa[9] ),
    .A(_04651_),
    .Y(_04786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1764 (.A(net1763),
    .X(net1764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10776_ (.Y(_04788_),
    .A(\fp16_res_pipe.add_renorm0.exp[5] ),
    .B(_04779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10777_ (.VDD(VPWR),
    .Y(_04789_),
    .A(_04788_),
    .VSS(VGND));
 sg13g2_nand2_1 _10778_ (.Y(_04790_),
    .A(_04786_),
    .B(\fp16_res_pipe.add_renorm0.exp[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10779_ (.B1(_04790_),
    .VDD(VPWR),
    .Y(_04791_),
    .VSS(VGND),
    .A1(_04786_),
    .A2(_04789_));
 sg13g2_buf_1 fanout130 (.A(net131),
    .X(net130),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10781_ (.Y(_04793_),
    .A(_03580_),
    .B(_04778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10782_ (.VDD(VPWR),
    .Y(_04794_),
    .A(_04793_),
    .VSS(VGND));
 sg13g2_nor2_1 _10783_ (.A(\fp16_res_pipe.add_renorm0.exp[4] ),
    .B(net1709),
    .Y(_04795_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _10784_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_04795_),
    .Y(_04796_),
    .A2(_04794_),
    .A1(net1709));
 sg13g2_nor2_1 _10785_ (.A(_04791_),
    .B(_04796_),
    .Y(_04797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10786_ (.VDD(VPWR),
    .Y(_04798_),
    .A(_04797_),
    .VSS(VGND));
 sg13g2_xnor2_1 _10787_ (.Y(_04799_),
    .A(\fp16_res_pipe.add_renorm0.exp[3] ),
    .B(_04777_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10788_ (.VDD(VPWR),
    .Y(_04800_),
    .A(_04799_),
    .VSS(VGND));
 sg13g2_nor2_1 _10789_ (.A(\fp16_res_pipe.add_renorm0.exp[3] ),
    .B(net1709),
    .Y(_04801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _10790_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_04801_),
    .Y(_04802_),
    .A2(_04800_),
    .A1(net1709));
 sg13g2_inv_1 _10791_ (.VDD(VPWR),
    .Y(_04803_),
    .A(\fp16_res_pipe.add_renorm0.exp[0] ),
    .VSS(VGND));
 sg13g2_o21ai_1 _10792_ (.B1(_03584_),
    .VDD(VPWR),
    .Y(_04804_),
    .VSS(VGND),
    .A1(_03586_),
    .A2(_04803_));
 sg13g2_and2_1 _10793_ (.A(_04804_),
    .B(_04777_),
    .X(_04805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10794_ (.VDD(VPWR),
    .Y(_04806_),
    .A(_04805_),
    .VSS(VGND));
 sg13g2_nor2_1 _10795_ (.A(\fp16_res_pipe.add_renorm0.exp[2] ),
    .B(_04775_),
    .Y(_04807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _10796_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_04807_),
    .Y(_04808_),
    .A2(_04806_),
    .A1(_04775_));
 sg13g2_inv_2 _10797_ (.Y(_04809_),
    .A(_04808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10798_ (.Y(_04810_),
    .A(_04809_),
    .B(_04740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10799_ (.A(_04802_),
    .B(_04810_),
    .Y(_04811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10800_ (.VDD(VPWR),
    .Y(_04812_),
    .A(_04811_),
    .VSS(VGND));
 sg13g2_nor2_1 _10801_ (.A(_04798_),
    .B(_04812_),
    .Y(_04813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10802_ (.Y(_04814_),
    .A(_03576_),
    .B(_04780_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10803_ (.VDD(VPWR),
    .Y(_04815_),
    .A(_04814_),
    .VSS(VGND));
 sg13g2_nor2_1 _10804_ (.A(\fp16_res_pipe.add_renorm0.exp[6] ),
    .B(net1709),
    .Y(_04816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _10805_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_04816_),
    .Y(_04817_),
    .A2(_04815_),
    .A1(net1709));
 sg13g2_inv_1 _10806_ (.VDD(VPWR),
    .Y(_04818_),
    .A(_04817_),
    .VSS(VGND));
 sg13g2_nand2_1 _10807_ (.Y(_04819_),
    .A(_04813_),
    .B(_04818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10808_ (.Y(_04820_),
    .A(_04785_),
    .B(_04819_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10809_ (.A(_04774_),
    .B(_04820_),
    .Y(_04821_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10810_ (.Y(_04822_),
    .A(_04809_),
    .B(_04724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10811_ (.Y(_04823_),
    .A(_04775_),
    .B(\fp16_res_pipe.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10812_ (.Y(_04824_),
    .A(\fp16_res_pipe.add_renorm0.exp[1] ),
    .B(_04823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10813_ (.A(_04822_),
    .B(_04824_),
    .X(_04825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04724_),
    .A2(_04808_),
    .Y(_04826_),
    .B1(_04825_));
 sg13g2_nor2_1 _10815_ (.A(_04796_),
    .B(_04802_),
    .Y(_04827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10816_ (.Y(_04828_),
    .A(_04826_),
    .B(_04827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10817_ (.VDD(VPWR),
    .Y(_04829_),
    .A(_04828_),
    .VSS(VGND));
 sg13g2_nor2_1 _10818_ (.A(_04791_),
    .B(_04817_),
    .Y(_04830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10819_ (.Y(_04831_),
    .A(_04829_),
    .B(_04830_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10820_ (.B1(_04743_),
    .VDD(VPWR),
    .Y(_04832_),
    .VSS(VGND),
    .A1(_04785_),
    .A2(_04831_));
 sg13g2_a21oi_1 _10821_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04831_),
    .A2(_04785_),
    .Y(_04833_),
    .B1(_04832_));
 sg13g2_nor3_1 _10822_ (.A(net1772),
    .B(_04821_),
    .C(_04833_),
    .Y(_04834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10823_ (.Y(_04835_),
    .A(_04809_),
    .B(_04735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10824_ (.VDD(VPWR),
    .Y(_04836_),
    .A(_04835_),
    .VSS(VGND));
 sg13g2_inv_2 _10825_ (.Y(_04837_),
    .A(_04824_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10826_ (.Y(_04838_),
    .A(_04722_),
    .B(_04734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10827_ (.Y(_04839_),
    .A(_04838_),
    .B(_04667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10828_ (.A(_04837_),
    .B(_04839_),
    .Y(_04840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10829_ (.Y(_04841_),
    .A(\fp16_res_pipe.add_renorm0.exp[0] ),
    .B(_04786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10830_ (.VDD(VPWR),
    .Y(_04842_),
    .A(_04841_),
    .VSS(VGND));
 sg13g2_xnor2_1 _10831_ (.Y(_04843_),
    .A(_04837_),
    .B(_04839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10832_ (.A(_04842_),
    .B(_04843_),
    .Y(_04844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10833_ (.A(_04840_),
    .B(_04844_),
    .Y(_04845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10834_ (.A(_04836_),
    .B(_04845_),
    .Y(_04846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10835_ (.Y(_04847_),
    .A(_04735_),
    .B(_04808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _10836_ (.A(_04846_),
    .B_N(_04847_),
    .Y(_04848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10837_ (.Y(_04849_),
    .A(_04802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _10838_ (.Y(_04850_),
    .A(_04848_),
    .B(_04849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _10839_ (.A(_04798_),
    .B(_04850_),
    .Y(_04851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10840_ (.VDD(VPWR),
    .Y(_04852_),
    .A(_04851_),
    .VSS(VGND));
 sg13g2_o21ai_1 _10841_ (.B1(_04785_),
    .VDD(VPWR),
    .Y(_04853_),
    .VSS(VGND),
    .A1(_04817_),
    .A2(_04852_));
 sg13g2_nand3_1 _10842_ (.B(_04784_),
    .C(_04818_),
    .A(_04851_),
    .Y(_04854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10843_ (.B(_04854_),
    .C(_04737_),
    .A(_04853_),
    .Y(_04855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10844_ (.Y(_04856_),
    .A(_04834_),
    .B(_04855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10845_ (.A(net1825),
    .B(\fp16_res_pipe.add_renorm0.exp[7] ),
    .Y(_04857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04782_),
    .A2(net1825),
    .Y(_04858_),
    .B1(_04857_));
 sg13g2_nor2_1 _10847_ (.A(net1825),
    .B(_03576_),
    .Y(_04859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04814_),
    .A2(net1825),
    .Y(_04860_),
    .B1(_04859_));
 sg13g2_nor2_1 _10849_ (.A(net1825),
    .B(_03580_),
    .Y(_04861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04793_),
    .A2(net1825),
    .Y(_04862_),
    .B1(_04861_));
 sg13g2_nor2_1 _10851_ (.A(net1824),
    .B(\fp16_res_pipe.add_renorm0.exp[0] ),
    .Y(_04863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10852_ (.Y(_04864_),
    .A(net1824),
    .B(\fp16_res_pipe.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _10853_ (.A(_04863_),
    .B_N(_04864_),
    .Y(_04865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10854_ (.Y(_04866_),
    .A(_04748_),
    .B(_04865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10855_ (.A(_03586_),
    .B(_04866_),
    .Y(_04867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10856_ (.A(net1824),
    .B(\fp16_res_pipe.add_renorm0.exp[2] ),
    .Y(_04868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10857_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04806_),
    .A2(net1824),
    .Y(_04869_),
    .B1(_04868_));
 sg13g2_nand2_1 _10858_ (.Y(_04870_),
    .A(_04867_),
    .B(_04869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10859_ (.VDD(VPWR),
    .Y(_04871_),
    .A(_04870_),
    .VSS(VGND));
 sg13g2_nor2_1 _10860_ (.A(net1824),
    .B(\fp16_res_pipe.add_renorm0.exp[3] ),
    .Y(_04872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10861_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04800_),
    .A2(net1824),
    .Y(_04873_),
    .B1(_04872_));
 sg13g2_nand2_1 _10862_ (.Y(_04874_),
    .A(_04871_),
    .B(_04873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10863_ (.A(_04862_),
    .B(_04874_),
    .Y(_04875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10864_ (.A(net1825),
    .B(\fp16_res_pipe.add_renorm0.exp[5] ),
    .Y(_04876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10865_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04789_),
    .A2(net1825),
    .Y(_04877_),
    .B1(_04876_));
 sg13g2_nand2_1 _10866_ (.Y(_04878_),
    .A(_04875_),
    .B(_04877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10867_ (.A(_04860_),
    .B(_04878_),
    .Y(_04879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10868_ (.Y(_04880_),
    .A(_04858_),
    .B(_04879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10869_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1772),
    .A2(_04880_),
    .Y(_04881_),
    .B1(_04771_));
 sg13g2_nand2_1 _10870_ (.Y(_04882_),
    .A(_04856_),
    .B(_04881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10871_ (.Y(_04883_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10872_ (.Y(_01135_),
    .A(_04882_),
    .B(_04883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10873_ (.VDD(VPWR),
    .Y(_04884_),
    .A(_04813_),
    .VSS(VGND));
 sg13g2_nand2_1 _10874_ (.Y(_04885_),
    .A(_04884_),
    .B(_04817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10875_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04885_),
    .A2(_04819_),
    .Y(_04886_),
    .B1(_04774_));
 sg13g2_nand2_1 _10876_ (.Y(_04887_),
    .A(_04826_),
    .B(_04849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10877_ (.VDD(VPWR),
    .Y(_04888_),
    .A(_04887_),
    .VSS(VGND));
 sg13g2_nand2_1 _10878_ (.Y(_04889_),
    .A(_04888_),
    .B(_04797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10879_ (.Y(_04890_),
    .A(_04889_),
    .B(_04817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10880_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04890_),
    .A2(_04831_),
    .Y(_04891_),
    .B1(_04742_));
 sg13g2_nor3_1 _10881_ (.A(net1772),
    .B(_04886_),
    .C(_04891_),
    .Y(_04892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10882_ (.Y(_04893_),
    .A(_04852_),
    .B(_04818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10883_ (.Y(_04894_),
    .A(_04851_),
    .B(_04817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10884_ (.B(_04737_),
    .C(_04894_),
    .A(_04893_),
    .Y(_04895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10885_ (.Y(_04896_),
    .A(_04892_),
    .B(_04895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _10886_ (.Y(_04897_),
    .A(_04771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10887_ (.A(_04878_),
    .B(_04860_),
    .X(_04898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10888_ (.B1(net1772),
    .VDD(VPWR),
    .Y(_04899_),
    .VSS(VGND),
    .A1(_04879_),
    .A2(_04898_));
 sg13g2_nand3_1 _10889_ (.B(_04897_),
    .C(_04899_),
    .A(_04896_),
    .Y(_04900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10890_ (.Y(_04901_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10891_ (.Y(_01134_),
    .A(_04900_),
    .B(_04901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10892_ (.VDD(VPWR),
    .Y(_04902_),
    .A(\fp16_res_pipe.y[12] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10893_ (.A(_04796_),
    .B(_04850_),
    .Y(_04903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _10894_ (.A(_04903_),
    .B_N(_04791_),
    .Y(_04904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10895_ (.B1(_04737_),
    .VDD(VPWR),
    .Y(_04905_),
    .VSS(VGND),
    .A1(_04851_),
    .A2(_04904_));
 sg13g2_o21ai_1 _10896_ (.B1(_04791_),
    .VDD(VPWR),
    .Y(_04906_),
    .VSS(VGND),
    .A1(_04796_),
    .A2(_04812_));
 sg13g2_a21oi_1 _10897_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04906_),
    .A2(_04884_),
    .Y(_04907_),
    .B1(_04774_));
 sg13g2_nand2_1 _10898_ (.Y(_04908_),
    .A(_04828_),
    .B(_04791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10899_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04889_),
    .A2(_04908_),
    .Y(_04909_),
    .B1(_04742_));
 sg13g2_nor3_1 _10900_ (.A(net1772),
    .B(_04907_),
    .C(_04909_),
    .Y(_04910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10901_ (.Y(_04911_),
    .A(_04905_),
    .B(_04910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _10902_ (.Y(_04912_),
    .A(_04877_),
    .B(_04875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10903_ (.Y(_04913_),
    .A(_04912_),
    .B(net1772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10904_ (.B(_04897_),
    .C(_04913_),
    .A(_04911_),
    .Y(_04914_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10905_ (.B1(_04914_),
    .VDD(VPWR),
    .Y(_01133_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.reg3en.q[0] ),
    .A2(_04902_));
 sg13g2_inv_1 _10906_ (.VDD(VPWR),
    .Y(_04915_),
    .A(_04796_),
    .VSS(VGND));
 sg13g2_inv_1 _10907_ (.VDD(VPWR),
    .Y(_04916_),
    .A(_04850_),
    .VSS(VGND));
 sg13g2_nor2_1 _10908_ (.A(_04915_),
    .B(_04916_),
    .Y(_04917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10909_ (.B1(_04737_),
    .VDD(VPWR),
    .Y(_04918_),
    .VSS(VGND),
    .A1(_04903_),
    .A2(_04917_));
 sg13g2_xnor2_1 _10910_ (.Y(_04919_),
    .A(_04915_),
    .B(_04811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10911_ (.Y(_04920_),
    .A(_04919_),
    .B(_04741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10912_ (.A(_04915_),
    .B(_04888_),
    .Y(_04921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10913_ (.B1(_04743_),
    .VDD(VPWR),
    .Y(_04922_),
    .VSS(VGND),
    .A1(_04829_),
    .A2(_04921_));
 sg13g2_nand4_1 _10914_ (.B(net1821),
    .C(_04920_),
    .A(_04918_),
    .Y(_04923_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04922_));
 sg13g2_inv_1 _10915_ (.VDD(VPWR),
    .Y(_04924_),
    .A(_04874_),
    .VSS(VGND));
 sg13g2_nor2b_1 _10916_ (.A(_04924_),
    .B_N(_04862_),
    .Y(_04925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10917_ (.B1(net1771),
    .VDD(VPWR),
    .Y(_04926_),
    .VSS(VGND),
    .A1(_04875_),
    .A2(_04925_));
 sg13g2_nand3_1 _10918_ (.B(_04897_),
    .C(_04926_),
    .A(_04923_),
    .Y(_04927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10919_ (.Y(_04928_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10920_ (.Y(_01132_),
    .A(_04927_),
    .B(_04928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _10921_ (.VDD(VPWR),
    .Y(_04929_),
    .A(\fp16_res_pipe.y[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _10922_ (.A(_04849_),
    .B(_04848_),
    .Y(_04930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10923_ (.B1(_04737_),
    .VDD(VPWR),
    .Y(_04931_),
    .VSS(VGND),
    .A1(_04930_),
    .A2(_04916_));
 sg13g2_a21oi_1 _10924_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04809_),
    .A2(_04740_),
    .Y(_04932_),
    .B1(_04849_));
 sg13g2_o21ai_1 _10925_ (.B1(_04741_),
    .VDD(VPWR),
    .Y(_04933_),
    .VSS(VGND),
    .A1(_04811_),
    .A2(_04932_));
 sg13g2_nor2_1 _10926_ (.A(_04849_),
    .B(_04826_),
    .Y(_04934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10927_ (.B1(_04743_),
    .VDD(VPWR),
    .Y(_04935_),
    .VSS(VGND),
    .A1(_04934_),
    .A2(_04888_));
 sg13g2_nand4_1 _10928_ (.B(net1821),
    .C(_04933_),
    .A(_04931_),
    .Y(_04936_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04935_));
 sg13g2_nor2_1 _10929_ (.A(_04873_),
    .B(_04871_),
    .Y(_04937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10930_ (.B1(net1771),
    .VDD(VPWR),
    .Y(_04938_),
    .VSS(VGND),
    .A1(_04937_),
    .A2(_04924_));
 sg13g2_nand3_1 _10931_ (.B(_04897_),
    .C(_04938_),
    .A(_04936_),
    .Y(_04939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10932_ (.B1(_04939_),
    .VDD(VPWR),
    .Y(_01131_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.reg3en.q[0] ),
    .A2(_04929_));
 sg13g2_inv_1 _10933_ (.VDD(VPWR),
    .Y(_04940_),
    .A(\fp16_res_pipe.y[9] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _10934_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04845_),
    .A2(_04836_),
    .Y(_04941_),
    .B1(_04739_));
 sg13g2_nand2b_1 _10935_ (.Y(_04942_),
    .B(_04941_),
    .A_N(_04846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10936_ (.A(_04740_),
    .B(_04809_),
    .Y(_04943_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10937_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04694_),
    .A2(_04809_),
    .Y(_04944_),
    .B1(_04943_));
 sg13g2_nor2_1 _10938_ (.A(_04742_),
    .B(_04825_),
    .Y(_04945_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10939_ (.B1(_04945_),
    .VDD(VPWR),
    .Y(_04946_),
    .VSS(VGND),
    .A1(_04824_),
    .A2(_04822_));
 sg13g2_nand4_1 _10940_ (.B(net1821),
    .C(_04944_),
    .A(_04942_),
    .Y(_04947_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_04946_));
 sg13g2_nor2_1 _10941_ (.A(_04869_),
    .B(_04867_),
    .Y(_04948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10942_ (.B1(net1771),
    .VDD(VPWR),
    .Y(_04949_),
    .VSS(VGND),
    .A1(_04948_),
    .A2(_04871_));
 sg13g2_nand3_1 _10943_ (.B(_04947_),
    .C(_04949_),
    .A(_04897_),
    .Y(_04950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10944_ (.B1(_04950_),
    .VDD(VPWR),
    .Y(_01130_),
    .VSS(VGND),
    .A1(\fp16_res_pipe.reg3en.q[0] ),
    .A2(_04940_));
 sg13g2_nand2_1 _10945_ (.Y(_04951_),
    .A(_04843_),
    .B(_04842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _10946_ (.B(_04737_),
    .C(_04951_),
    .Y(_04952_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_04844_));
 sg13g2_o21ai_1 _10947_ (.B1(\fp16_res_pipe.seg_reg1.q[21] ),
    .VDD(VPWR),
    .Y(_04953_),
    .VSS(VGND),
    .A1(_04837_),
    .A2(_04774_));
 sg13g2_a21oi_1 _10948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04743_),
    .A2(_04837_),
    .Y(_04954_),
    .B1(_04953_));
 sg13g2_inv_1 _10949_ (.VDD(VPWR),
    .Y(_04955_),
    .A(_04748_),
    .VSS(VGND));
 sg13g2_a21oi_1 _10950_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04955_),
    .A2(_04864_),
    .Y(_04956_),
    .B1(_04863_));
 sg13g2_nor2_1 _10951_ (.A(_03586_),
    .B(_04956_),
    .Y(_04957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _10952_ (.A(_04956_),
    .B(_03586_),
    .X(_04958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _10953_ (.A(\fp16_res_pipe.seg_reg1.q[21] ),
    .B(_04957_),
    .C(_04958_),
    .Y(_04959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _10954_ (.A2(_04954_),
    .A1(_04952_),
    .B1(_04959_),
    .X(_04960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10955_ (.Y(_04961_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10956_ (.B1(_04961_),
    .VDD(VPWR),
    .Y(_01129_),
    .VSS(VGND),
    .A1(_04960_),
    .A2(_04771_));
 sg13g2_nand2b_1 _10957_ (.Y(_04962_),
    .B(_04955_),
    .A_N(_04865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10958_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04748_),
    .A2(_04865_),
    .Y(_04963_),
    .B1(\fp16_res_pipe.seg_reg1.q[21] ));
 sg13g2_nand2_1 _10959_ (.Y(_04964_),
    .A(_04739_),
    .B(_04842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10960_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04744_),
    .A2(_04841_),
    .Y(_04965_),
    .B1(net1771));
 sg13g2_a22oi_1 _10961_ (.Y(_04966_),
    .B1(_04964_),
    .B2(_04965_),
    .A2(_04963_),
    .A1(_04962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10962_ (.Y(_04967_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10963_ (.B1(_04967_),
    .VDD(VPWR),
    .Y(_01128_),
    .VSS(VGND),
    .A1(_04966_),
    .A2(_04771_));
 sg13g2_mux2_1 _10964_ (.A0(\fp16_res_pipe.y[6] ),
    .A1(_04732_),
    .S(net1835),
    .X(_01127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _10965_ (.A0(\fp16_res_pipe.y[5] ),
    .A1(_04768_),
    .S(\fp16_res_pipe.reg3en.q[0] ),
    .X(_01126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _10966_ (.A0(\fp16_res_pipe.y[4] ),
    .A1(_04702_),
    .S(net1835),
    .X(_01125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _10967_ (.A0(\fp16_res_pipe.y[3] ),
    .A1(_04686_),
    .S(net1835),
    .X(_01124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10968_ (.Y(_04968_),
    .A(_04670_),
    .B(_04695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10969_ (.Y(_04969_),
    .A(_04679_),
    .B(_04672_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10970_ (.Y(_04970_),
    .A(net1710),
    .B(_04681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _10971_ (.B(_04969_),
    .C(_04970_),
    .A(_04968_),
    .Y(_04971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _10972_ (.A(net1821),
    .B(_04756_),
    .Y(_04972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10973_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04971_),
    .A2(net1821),
    .Y(_04973_),
    .B1(_04972_));
 sg13g2_nor2_1 _10974_ (.A(net1835),
    .B(\fp16_res_pipe.y[2] ),
    .Y(_04974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _10975_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04973_),
    .A2(net1835),
    .Y(_01123_),
    .B1(_04974_));
 sg13g2_mux2_1 _10976_ (.A0(\fp16_res_pipe.y[1] ),
    .A1(_04708_),
    .S(net1835),
    .X(_01122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10977_ (.Y(_04975_),
    .A(_04772_),
    .B(\fp16_res_pipe.y[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10978_ (.B1(_04975_),
    .VDD(VPWR),
    .Y(_01121_),
    .VSS(VGND),
    .A1(_04772_),
    .A2(_04759_));
 sg13g2_mux2_1 _10979_ (.A0(\fp16_sum_pipe.exp_mant_logic0.b[15] ),
    .A1(\fp16_res_pipe.x2[15] ),
    .S(net1930),
    .X(_01120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _10980_ (.Y(_04976_),
    .A(\fp16_res_pipe.x2[14] ),
    .B(net1926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10981_ (.B1(_04976_),
    .VDD(VPWR),
    .Y(_01119_),
    .VSS(VGND),
    .A1(net1926),
    .A2(_02463_));
 sg13g2_nand2_1 _10982_ (.Y(_04977_),
    .A(\fp16_res_pipe.x2[13] ),
    .B(net1925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10983_ (.B1(_04977_),
    .VDD(VPWR),
    .Y(_01118_),
    .VSS(VGND),
    .A1(net1925),
    .A2(_02464_));
 sg13g2_nand2_1 _10984_ (.Y(_04978_),
    .A(\fp16_res_pipe.x2[12] ),
    .B(net1924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10985_ (.B1(_04978_),
    .VDD(VPWR),
    .Y(_01117_),
    .VSS(VGND),
    .A1(net1926),
    .A2(_02199_));
 sg13g2_nand2_1 _10986_ (.Y(_04979_),
    .A(\fp16_res_pipe.x2[11] ),
    .B(net1924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10987_ (.B1(_04979_),
    .VDD(VPWR),
    .Y(_01116_),
    .VSS(VGND),
    .A1(net1926),
    .A2(_02194_));
 sg13g2_nand2_1 _10988_ (.Y(_04980_),
    .A(\fp16_res_pipe.x2[10] ),
    .B(net1931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10989_ (.B1(_04980_),
    .VDD(VPWR),
    .Y(_01115_),
    .VSS(VGND),
    .A1(net1931),
    .A2(_02205_));
 sg13g2_nand2_1 _10990_ (.Y(_04981_),
    .A(\fp16_res_pipe.x2[9] ),
    .B(net1932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10991_ (.B1(_04981_),
    .VDD(VPWR),
    .Y(_01114_),
    .VSS(VGND),
    .A1(net1933),
    .A2(_02210_));
 sg13g2_nand2_1 _10992_ (.Y(_04982_),
    .A(\fp16_res_pipe.x2[8] ),
    .B(net1932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10993_ (.B1(_04982_),
    .VDD(VPWR),
    .Y(_01113_),
    .VSS(VGND),
    .A1(net1932),
    .A2(_02227_));
 sg13g2_nand2_1 _10994_ (.Y(_04983_),
    .A(\fp16_res_pipe.x2[7] ),
    .B(net1933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10995_ (.B1(_04983_),
    .VDD(VPWR),
    .Y(_01112_),
    .VSS(VGND),
    .A1(net1933),
    .A2(_02216_));
 sg13g2_nand2_1 _10996_ (.Y(_04984_),
    .A(\fp16_res_pipe.x2[6] ),
    .B(net1928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10997_ (.B1(_04984_),
    .VDD(VPWR),
    .Y(_01111_),
    .VSS(VGND),
    .A1(net1929),
    .A2(_02466_));
 sg13g2_nand2_1 _10998_ (.Y(_04985_),
    .A(\fp16_res_pipe.x2[5] ),
    .B(net1927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _10999_ (.B1(_04985_),
    .VDD(VPWR),
    .Y(_01110_),
    .VSS(VGND),
    .A1(net1928),
    .A2(_02458_));
 sg13g2_nand2_1 _11000_ (.Y(_04986_),
    .A(\fp16_res_pipe.x2[4] ),
    .B(net1928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11001_ (.B1(_04986_),
    .VDD(VPWR),
    .Y(_01109_),
    .VSS(VGND),
    .A1(net1929),
    .A2(_02459_));
 sg13g2_nand2_1 _11002_ (.Y(_04987_),
    .A(\fp16_res_pipe.x2[3] ),
    .B(net1928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11003_ (.B1(_04987_),
    .VDD(VPWR),
    .Y(_01108_),
    .VSS(VGND),
    .A1(net1929),
    .A2(_02467_));
 sg13g2_nand2_1 _11004_ (.Y(_04988_),
    .A(\fp16_res_pipe.x2[2] ),
    .B(net1927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11005_ (.B1(_04988_),
    .VDD(VPWR),
    .Y(_01107_),
    .VSS(VGND),
    .A1(net1929),
    .A2(_02468_));
 sg13g2_nand2_1 _11006_ (.Y(_04989_),
    .A(\fp16_res_pipe.x2[1] ),
    .B(net1925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11007_ (.B1(_04989_),
    .VDD(VPWR),
    .Y(_01106_),
    .VSS(VGND),
    .A1(net1928),
    .A2(_02460_));
 sg13g2_nand2_1 _11008_ (.Y(_04990_),
    .A(\fp16_res_pipe.x2[0] ),
    .B(net1929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11009_ (.B1(_04990_),
    .VDD(VPWR),
    .Y(_01105_),
    .VSS(VGND),
    .A1(net1929),
    .A2(_02469_));
 sg13g2_nand2_1 _11010_ (.Y(_04991_),
    .A(\acc_sum.exp_mant_logic0.a[15] ),
    .B(net1813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11011_ (.B1(_04991_),
    .VDD(VPWR),
    .Y(_01104_),
    .VSS(VGND),
    .A1(net1813),
    .A2(_02802_));
 sg13g2_mux2_1 _11012_ (.A0(\acc_sum.op_sign_logic0.s_b ),
    .A1(\acc_sum.exp_mant_logic0.b[15] ),
    .S(net1813),
    .X(_01103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11013_ (.VDD(VPWR),
    .Y(_04992_),
    .A(\acc_sum.seg_reg0.q[29] ),
    .VSS(VGND));
 sg13g2_inv_4 _11014_ (.A(\acc_sum.reg1en.q[0] ),
    .Y(_04993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout59 (.A(net60),
    .X(net59),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout58 (.A(net60),
    .X(net58),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11017_ (.A(\acc_sum.exp_mant_logic0.b[14] ),
    .B(_04993_),
    .Y(_04996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11018_ (.Y(_04997_),
    .A(\acc_sum.exp_mant_logic0.a[14] ),
    .B(\acc_sum.exp_mant_logic0.b[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11019_ (.Y(_04998_),
    .A(_04997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11020_ (.A(\acc_sum.exp_mant_logic0.b[12] ),
    .B(_02939_),
    .Y(_04999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11021_ (.A(\acc_sum.exp_mant_logic0.a[12] ),
    .B(_03333_),
    .Y(_05000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11022_ (.A(_04999_),
    .B(_05000_),
    .Y(_05001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11023_ (.VDD(VPWR),
    .Y(_05002_),
    .A(_05001_),
    .VSS(VGND));
 sg13g2_nor2_1 _11024_ (.A(\acc_sum.exp_mant_logic0.b[11] ),
    .B(_02941_),
    .Y(_05003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11025_ (.A(\acc_sum.exp_mant_logic0.a[11] ),
    .B(_03335_),
    .Y(_05004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11026_ (.A(_05003_),
    .B(_05004_),
    .Y(_05005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11027_ (.VDD(VPWR),
    .Y(_05006_),
    .A(_05005_),
    .VSS(VGND));
 sg13g2_nor2_1 _11028_ (.A(\acc_sum.exp_mant_logic0.a[13] ),
    .B(_03331_),
    .Y(_05007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11029_ (.A(\acc_sum.exp_mant_logic0.b[13] ),
    .B(_02937_),
    .Y(_05008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11030_ (.Y(_05009_),
    .A(_05008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _11031_ (.Y(_05010_),
    .B(_05009_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05007_));
 sg13g2_nor4_1 _11032_ (.A(_04998_),
    .B(_05002_),
    .C(_05006_),
    .D(_05010_),
    .Y(_05011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11033_ (.A(\acc_sum.exp_mant_logic0.b[10] ),
    .B(_02943_),
    .Y(_05012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11034_ (.A(\acc_sum.exp_mant_logic0.a[10] ),
    .B(_03337_),
    .Y(_05013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11035_ (.A(_05012_),
    .B(_05013_),
    .Y(_05014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11036_ (.A(\acc_sum.exp_mant_logic0.b[9] ),
    .B(_02945_),
    .Y(_05015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11037_ (.A(\acc_sum.exp_mant_logic0.a[9] ),
    .B(_03339_),
    .Y(_05016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11038_ (.A(_05015_),
    .B(_05016_),
    .Y(_05017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11039_ (.Y(_05018_),
    .A(_05014_),
    .B(_05017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _11040_ (.B(\acc_sum.exp_mant_logic0.b[8] ),
    .A(\acc_sum.exp_mant_logic0.a[8] ),
    .X(_05019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11041_ (.VDD(VPWR),
    .Y(_05020_),
    .A(_05019_),
    .VSS(VGND));
 sg13g2_nor2_2 _11042_ (.A(\acc_sum.exp_mant_logic0.a[7] ),
    .B(_03343_),
    .Y(_05021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11043_ (.A(\acc_sum.exp_mant_logic0.b[7] ),
    .B(_02949_),
    .Y(_05022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11044_ (.A(_05021_),
    .B(_05022_),
    .Y(_05023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _11045_ (.Y(_05024_),
    .A(_05020_),
    .B(_05023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11046_ (.A(_05018_),
    .B(_05024_),
    .Y(_05025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _11047_ (.Y(_05026_),
    .A(_05011_),
    .B(_05025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1722 (.A(_07076_),
    .X(net1722),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11049_ (.Y(_05028_),
    .A(_05026_),
    .B(\acc_sum.exp_mant_logic0.a[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11050_ (.Y(_01102_),
    .B1(_04996_),
    .B2(_05028_),
    .A2(net1760),
    .A1(_04992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11051_ (.Y(_05029_),
    .A(_03341_),
    .B(\acc_sum.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11052_ (.B1(_05029_),
    .VDD(VPWR),
    .Y(_05030_),
    .VSS(VGND),
    .A1(_05021_),
    .A2(_05019_));
 sg13g2_inv_1 _11053_ (.VDD(VPWR),
    .Y(_05031_),
    .A(_05016_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11054_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05030_),
    .A2(_05031_),
    .Y(_05032_),
    .B1(_05015_));
 sg13g2_inv_1 _11055_ (.VDD(VPWR),
    .Y(_05033_),
    .A(_05012_),
    .VSS(VGND));
 sg13g2_o21ai_1 _11056_ (.B1(_05033_),
    .VDD(VPWR),
    .Y(_05034_),
    .VSS(VGND),
    .A1(_05013_),
    .A2(_05032_));
 sg13g2_nand2_1 _11057_ (.Y(_05035_),
    .A(_05034_),
    .B(_05011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11058_ (.A(_04998_),
    .B(_05010_),
    .Y(_05036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11059_ (.VDD(VPWR),
    .Y(_05037_),
    .A(_05003_),
    .VSS(VGND));
 sg13g2_inv_1 _11060_ (.VDD(VPWR),
    .Y(_05038_),
    .A(_04999_),
    .VSS(VGND));
 sg13g2_o21ai_1 _11061_ (.B1(_05038_),
    .VDD(VPWR),
    .Y(_05039_),
    .VSS(VGND),
    .A1(_05000_),
    .A2(_05037_));
 sg13g2_nor2_1 _11062_ (.A(_05009_),
    .B(_04998_),
    .Y(_05040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _11063_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_05039_),
    .C1(_05040_),
    .B1(_05036_),
    .A1(\acc_sum.exp_mant_logic0.a[14] ),
    .Y(_05041_),
    .A2(_03329_));
 sg13g2_nand2_2 _11064_ (.Y(_05042_),
    .A(_05035_),
    .B(_05041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout57 (.A(net60),
    .X(net57),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11066_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05042_),
    .A2(_02937_),
    .Y(_05044_),
    .B1(_04993_));
 sg13g2_o21ai_1 _11067_ (.B1(_05044_),
    .VDD(VPWR),
    .Y(_05045_),
    .VSS(VGND),
    .A1(\acc_sum.exp_mant_logic0.b[13] ),
    .A2(_05042_));
 sg13g2_o21ai_1 _11068_ (.B1(_05045_),
    .VDD(VPWR),
    .Y(_01101_),
    .VSS(VGND),
    .A1(_02922_),
    .A2(net1813));
 sg13g2_nand2_2 _11069_ (.Y(_05046_),
    .A(_05042_),
    .B(_05026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout133 (.A(net136),
    .X(net133),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11071_ (.Y(_05048_),
    .A(_05046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11072_ (.A(_04993_),
    .B(_05048_),
    .Y(_05049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _11073_ (.A(_05049_),
    .Y(_05050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout132 (.A(net136),
    .X(net132),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11075_ (.A(_04993_),
    .B(_05046_),
    .Y(_05052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11078_ (.Y(_05055_),
    .B1(\acc_sum.exp_mant_logic0.a[12] ),
    .B2(_05052_),
    .A2(_04993_),
    .A1(\acc_sum.seg_reg0.q[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11079_ (.B1(_05055_),
    .VDD(VPWR),
    .Y(_01100_),
    .VSS(VGND),
    .A1(_03333_),
    .A2(_05050_));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11081_ (.Y(_05057_),
    .A(_05049_),
    .B(\acc_sum.exp_mant_logic0.b[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11082_ (.Y(_05058_),
    .A(_05052_),
    .B(\acc_sum.exp_mant_logic0.a[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11083_ (.Y(_05059_),
    .A(_04993_),
    .B(\acc_sum.seg_reg0.q[26] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11084_ (.B(_05058_),
    .C(_05059_),
    .A(_05057_),
    .Y(_01099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11085_ (.Y(_05060_),
    .A(_05049_),
    .B(\acc_sum.exp_mant_logic0.b[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11086_ (.Y(_05061_),
    .A(_05052_),
    .B(\acc_sum.exp_mant_logic0.a[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11087_ (.Y(_05062_),
    .A(net1760),
    .B(\acc_sum.seg_reg0.q[25] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11088_ (.B(_05061_),
    .C(_05062_),
    .A(_05060_),
    .Y(_01098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11089_ (.Y(_05063_),
    .B1(\acc_sum.exp_mant_logic0.a[9] ),
    .B2(_05052_),
    .A2(net1760),
    .A1(\acc_sum.seg_reg0.q[24] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11090_ (.B1(_05063_),
    .VDD(VPWR),
    .Y(_01097_),
    .VSS(VGND),
    .A1(_03339_),
    .A2(_05050_));
 sg13g2_nand2_1 _11091_ (.Y(_05064_),
    .A(_05049_),
    .B(\acc_sum.exp_mant_logic0.b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11092_ (.Y(_05065_),
    .A(_05052_),
    .B(\acc_sum.exp_mant_logic0.a[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11093_ (.Y(_05066_),
    .A(net1760),
    .B(\acc_sum.seg_reg0.q[23] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11094_ (.B(_05065_),
    .C(_05066_),
    .A(_05064_),
    .Y(_01096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11095_ (.Y(_05067_),
    .B1(\acc_sum.exp_mant_logic0.a[7] ),
    .B2(_05052_),
    .A2(net1760),
    .A1(\acc_sum.seg_reg0.q[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11096_ (.B1(_05067_),
    .VDD(VPWR),
    .Y(_01095_),
    .VSS(VGND),
    .A1(_03343_),
    .A2(_05050_));
 sg13g2_nand3_1 _11097_ (.B(_02955_),
    .C(_02961_),
    .A(_02953_),
    .Y(_05068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11098_ (.B(_02945_),
    .C(_02947_),
    .A(_02943_),
    .Y(_05069_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02949_));
 sg13g2_nand4_1 _11099_ (.B(_02937_),
    .C(_02939_),
    .A(_02935_),
    .Y(_05070_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02941_));
 sg13g2_nand4_1 _11100_ (.B(_02957_),
    .C(_02959_),
    .A(_02951_),
    .Y(_05071_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02963_));
 sg13g2_nor4_2 _11101_ (.A(_05068_),
    .B(_05069_),
    .C(_05070_),
    .Y(_05072_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_05071_));
 sg13g2_inv_4 _11102_ (.A(_05072_),
    .Y(_05073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11103_ (.B(\acc_sum.reg1en.q[0] ),
    .C(_05073_),
    .A(_05042_),
    .Y(_05074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11104_ (.B1(_05074_),
    .VDD(VPWR),
    .Y(_01094_),
    .VSS(VGND),
    .A1(net1813),
    .A2(_02795_));
 sg13g2_inv_2 _11105_ (.Y(_05075_),
    .A(_05026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout134 (.A(net136),
    .X(net134),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11107_ (.Y(_05077_),
    .A(_02947_),
    .B(\acc_sum.exp_mant_logic0.b[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11108_ (.B1(_05077_),
    .VDD(VPWR),
    .Y(_05078_),
    .VSS(VGND),
    .A1(_05022_),
    .A2(_05019_));
 sg13g2_inv_1 _11109_ (.VDD(VPWR),
    .Y(_05079_),
    .A(_05078_),
    .VSS(VGND));
 sg13g2_nor2_1 _11110_ (.A(_05018_),
    .B(_05079_),
    .Y(_05080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11111_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05033_),
    .A2(_05016_),
    .Y(_05081_),
    .B1(_05013_));
 sg13g2_nor2b_1 _11112_ (.A(_05080_),
    .B_N(_05081_),
    .Y(_05082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11113_ (.VDD(VPWR),
    .Y(_05083_),
    .A(_05082_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05083_),
    .A2(_05005_),
    .Y(_05084_),
    .B1(_05004_));
 sg13g2_inv_1 _11115_ (.VDD(VPWR),
    .Y(_05085_),
    .A(_05084_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05085_),
    .A2(_05038_),
    .Y(_05086_),
    .B1(_05000_));
 sg13g2_inv_1 _11117_ (.VDD(VPWR),
    .Y(_05087_),
    .A(_05086_),
    .VSS(VGND));
 sg13g2_o21ai_1 _11118_ (.B1(_05009_),
    .VDD(VPWR),
    .Y(_05088_),
    .VSS(VGND),
    .A1(_05007_),
    .A2(_05087_));
 sg13g2_a21oi_1 _11119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05034_),
    .A2(_05005_),
    .Y(_05089_),
    .B1(_05003_));
 sg13g2_o21ai_1 _11120_ (.B1(_05038_),
    .VDD(VPWR),
    .Y(_05090_),
    .VSS(VGND),
    .A1(_05000_),
    .A2(_05089_));
 sg13g2_nand2b_1 _11121_ (.Y(_05091_),
    .B(_05090_),
    .A_N(_05007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11122_ (.Y(_05092_),
    .B1(_05009_),
    .B2(_05091_),
    .A2(\acc_sum.exp_mant_logic0.b[14] ),
    .A1(_02935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11123_ (.Y(_05093_),
    .A(_05092_),
    .B(_05026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11124_ (.B1(_05093_),
    .VDD(VPWR),
    .Y(_05094_),
    .VSS(VGND),
    .A1(_05048_),
    .A2(_05088_));
 sg13g2_nand2_1 _11125_ (.Y(_05095_),
    .A(_05094_),
    .B(_04998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11126_ (.A(_05034_),
    .B(net1698),
    .Y(_05096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05046_),
    .A2(_05082_),
    .Y(_05097_),
    .B1(_05096_));
 sg13g2_xnor2_1 _11128_ (.Y(_05098_),
    .A(_05006_),
    .B(_05097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11129_ (.Y(_05099_),
    .A(net1698),
    .B(_05085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11130_ (.B1(_05099_),
    .VDD(VPWR),
    .Y(_05100_),
    .VSS(VGND),
    .A1(_05089_),
    .A2(_05046_));
 sg13g2_xnor2_1 _11131_ (.Y(_05101_),
    .A(_05002_),
    .B(_05100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11132_ (.A(_05086_),
    .B(_05048_),
    .Y(_05102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11133_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05090_),
    .A2(_05048_),
    .Y(_05103_),
    .B1(_05102_));
 sg13g2_xor2_1 _11134_ (.B(_05103_),
    .A(_05010_),
    .X(_05104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11135_ (.A(_05098_),
    .B(_05101_),
    .C(_05104_),
    .Y(_05105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _11136_ (.Y(_05106_),
    .A(_05095_),
    .B(_05105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_49_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_49_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11138_ (.Y(_05108_),
    .B(net1698),
    .A_N(_05022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11139_ (.B1(_05108_),
    .VDD(VPWR),
    .Y(_05109_),
    .VSS(VGND),
    .A1(_05021_),
    .A2(net1698));
 sg13g2_xnor2_1 _11140_ (.Y(_05110_),
    .A(_05019_),
    .B(_05109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11141_ (.A(_05023_),
    .B(_05110_),
    .Y(_05111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11142_ (.Y(_05112_),
    .A(_05111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11143_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05079_),
    .A2(_05031_),
    .Y(_05113_),
    .B1(_05015_));
 sg13g2_nand2_1 _11144_ (.Y(_05114_),
    .A(net1698),
    .B(_05113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11145_ (.B1(_05114_),
    .VDD(VPWR),
    .Y(_05115_),
    .VSS(VGND),
    .A1(_05032_),
    .A2(net1698));
 sg13g2_xor2_1 _11146_ (.B(_05115_),
    .A(_05014_),
    .X(_05116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11147_ (.Y(_05117_),
    .A(net1698),
    .B(_05079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11148_ (.B1(_05117_),
    .VDD(VPWR),
    .Y(_05118_),
    .VSS(VGND),
    .A1(_05030_),
    .A2(net1698));
 sg13g2_xor2_1 _11149_ (.B(_05118_),
    .A(_05017_),
    .X(_05119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11150_ (.VDD(VPWR),
    .Y(_05120_),
    .A(_05119_),
    .VSS(VGND));
 sg13g2_nor2_1 _11151_ (.A(_05116_),
    .B(_05120_),
    .Y(_05121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11152_ (.Y(_05122_),
    .A(_05121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11153_ (.A(_05112_),
    .B(_05122_),
    .Y(_05123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11154_ (.A(net1663),
    .B_N(_05123_),
    .Y(_05124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_62_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_62_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11156_ (.Y(_05126_),
    .B1(_05073_),
    .B2(_05124_),
    .A2(_05075_),
    .A1(net1808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11157_ (.Y(_05127_),
    .B(_05046_),
    .A_N(_05126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11158_ (.Y(_05128_),
    .B1(net1808),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[9] ),
    .A1(net1760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11159_ (.B1(_05128_),
    .VDD(VPWR),
    .Y(_01093_),
    .VSS(VGND),
    .A1(net1760),
    .A2(_05127_));
 sg13g2_nor3_1 _11160_ (.A(_05024_),
    .B(_05120_),
    .C(_05106_),
    .Y(_05129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11161_ (.VDD(VPWR),
    .Y(_05130_),
    .A(_05106_),
    .VSS(VGND));
 sg13g2_nor2_1 _11162_ (.A(_05119_),
    .B(_05116_),
    .Y(_05131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11163_ (.B(_05024_),
    .C(_05131_),
    .A(_05130_),
    .Y(_05132_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11164_ (.Y(_05133_),
    .B(_05132_),
    .A_N(_05129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11165_ (.Y(_05134_),
    .A(_05023_),
    .B(_05019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11166_ (.A(_05134_),
    .B(_05122_),
    .Y(_05135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _11167_ (.A(net1663),
    .B_N(_05135_),
    .Y(_05136_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_67_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_67_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11169_ (.A(_05124_),
    .B(_05136_),
    .Y(_05138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11170_ (.Y(_05139_),
    .B(_05110_),
    .A_N(_05023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11171_ (.A(_05139_),
    .B(_05122_),
    .Y(_05140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11172_ (.A(net1663),
    .B_N(_05140_),
    .Y(_05141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_69_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_69_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11174_ (.Y(_05143_),
    .A(_05141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11175_ (.Y(_05144_),
    .A(_05131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11176_ (.A(_05024_),
    .B(_05144_),
    .Y(_05145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11177_ (.A(net1663),
    .B_N(_05145_),
    .Y(_05146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_51_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_51_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11179_ (.Y(_05148_),
    .A(_05146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11180_ (.B(_05143_),
    .C(_05148_),
    .A(_05138_),
    .Y(_05149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11181_ (.A(_05133_),
    .B(_05149_),
    .Y(_05150_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11182_ (.A(_05050_),
    .B(_05150_),
    .Y(_05151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_101_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_101_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_66_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_66_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11185_ (.Y(_05154_),
    .A(net1655),
    .B(_05073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11186_ (.Y(_05155_),
    .A(_05124_),
    .B(net1808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11187_ (.Y(_05156_),
    .A(_05075_),
    .B(net1809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11188_ (.B(_05155_),
    .C(_05156_),
    .A(_05154_),
    .Y(_05157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11189_ (.Y(_05158_),
    .A(net1635),
    .B(_05157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11190_ (.Y(_05159_),
    .B1(net1809),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[8] ),
    .A1(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11191_ (.Y(_01092_),
    .A(_05158_),
    .B(_05159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_68_clk (.A(clknet_5_28__leaf_clk),
    .X(clknet_leaf_68_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _11193_ (.A(_05122_),
    .B(_05112_),
    .C(net1663),
    .Y(_05161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11194_ (.Y(_05162_),
    .B1(net1809),
    .B2(_05161_),
    .A2(_05141_),
    .A1(_05073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11195_ (.Y(_05163_),
    .B1(net1808),
    .B2(net1655),
    .A2(_05075_),
    .A1(net1810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11196_ (.Y(_05164_),
    .A(_05162_),
    .B(_05163_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11197_ (.Y(_05165_),
    .A(net1635),
    .B(_05164_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11198_ (.Y(_05166_),
    .B1(net1810),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[7] ),
    .A1(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11199_ (.Y(_01091_),
    .A(_05165_),
    .B(_05166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11200_ (.Y(_05167_),
    .B1(_05073_),
    .B2(net1661),
    .A2(net1808),
    .A1(_05141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11201_ (.Y(_05168_),
    .B1(net1809),
    .B2(net1655),
    .A2(net1810),
    .A1(_05124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11202_ (.Y(_05169_),
    .A(_05075_),
    .B(\acc_sum.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11203_ (.B(_05168_),
    .C(_05169_),
    .A(_05167_),
    .Y(_05170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11204_ (.Y(_05171_),
    .A(net1635),
    .B(_05170_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11205_ (.Y(_05172_),
    .B1(\acc_sum.exp_mant_logic0.a[3] ),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[6] ),
    .A1(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11206_ (.Y(_01090_),
    .A(_05171_),
    .B(_05172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11207_ (.Y(_05173_),
    .A(net1655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11208_ (.A(_02955_),
    .B(_05173_),
    .Y(_05174_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11209_ (.A(_02951_),
    .B(_05148_),
    .Y(_05175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11210_ (.B(_05121_),
    .C(_05111_),
    .A(_05130_),
    .Y(_05176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11211_ (.A(_02957_),
    .B(_05176_),
    .Y(_05177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11212_ (.A(_05174_),
    .B(_05175_),
    .C(_05177_),
    .Y(_05178_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11213_ (.A(_02959_),
    .B(_05026_),
    .Y(_05179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11214_ (.A(_05112_),
    .B(_05144_),
    .Y(_05180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11215_ (.A(net1663),
    .B_N(_05180_),
    .Y(_05181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_70_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_70_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11217_ (.VDD(VPWR),
    .Y(_05183_),
    .A(_05181_),
    .VSS(VGND));
 sg13g2_nor2_1 _11218_ (.A(_05072_),
    .B(_05183_),
    .Y(_05184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11219_ (.A(_02953_),
    .B(_05143_),
    .Y(_05185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11220_ (.A(_05179_),
    .B(_05184_),
    .C(_05185_),
    .Y(_05186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11221_ (.Y(_05187_),
    .A(_05178_),
    .B(_05186_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11222_ (.Y(_05188_),
    .A(_05151_),
    .B(_05187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11223_ (.Y(_05189_),
    .B1(\acc_sum.exp_mant_logic0.a[2] ),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[5] ),
    .A1(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11224_ (.Y(_01089_),
    .A(_05188_),
    .B(_05189_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11225_ (.A(_02957_),
    .B(_05173_),
    .Y(_05190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11226_ (.A(_05134_),
    .B(_05144_),
    .Y(_05191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11227_ (.A(net1663),
    .B_N(_05191_),
    .Y(_05192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1658 (.A(_02347_),
    .X(net1658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11229_ (.Y(_05194_),
    .A(_05192_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11230_ (.A(_05072_),
    .B(_05194_),
    .Y(_05195_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11231_ (.A(_02953_),
    .B(_05148_),
    .Y(_05196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11232_ (.A(_05190_),
    .B(_05195_),
    .C(_05196_),
    .Y(_05197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11233_ (.Y(_05198_),
    .B1(\acc_sum.exp_mant_logic0.a[2] ),
    .B2(_05161_),
    .A2(net1653),
    .A1(net1808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11234_ (.Y(_05199_),
    .B1(net1810),
    .B2(_05141_),
    .A2(_05075_),
    .A1(\acc_sum.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11235_ (.B(_05198_),
    .C(_05199_),
    .A(_05197_),
    .Y(_05200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11236_ (.Y(_05201_),
    .A(_05200_),
    .B(net1635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11237_ (.Y(_05202_),
    .B1(\acc_sum.exp_mant_logic0.a[1] ),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[4] ),
    .A1(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11238_ (.Y(_01088_),
    .A(_05201_),
    .B(_05202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11239_ (.Y(_05203_),
    .A(net1661),
    .B(net1810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11240_ (.B1(_05203_),
    .VDD(VPWR),
    .Y(_05204_),
    .VSS(VGND),
    .A1(_02963_),
    .A2(_05026_));
 sg13g2_nand2_1 _11241_ (.Y(_05205_),
    .A(net1655),
    .B(\acc_sum.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11242_ (.B1(_05205_),
    .VDD(VPWR),
    .Y(_05206_),
    .VSS(VGND),
    .A1(_02957_),
    .A2(_05143_));
 sg13g2_nor2_1 _11243_ (.A(_05204_),
    .B(_05206_),
    .Y(_05207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11244_ (.Y(_05208_),
    .A(_05161_),
    .B(\acc_sum.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11245_ (.A(_02951_),
    .B(_05194_),
    .Y(_05209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11246_ (.A(_05139_),
    .B(_05144_),
    .Y(_05210_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11247_ (.A(net1663),
    .B_N(_05210_),
    .Y(_05211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_71_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_71_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11249_ (.Y(_05213_),
    .A(_05211_),
    .B(_05073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11250_ (.Y(_05214_),
    .A(net1653),
    .B(net1809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11251_ (.Y(_05215_),
    .A(_05213_),
    .B(_05214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11252_ (.A(_05209_),
    .B(_05215_),
    .Y(_05216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11253_ (.B(_05208_),
    .C(_05216_),
    .A(_05207_),
    .Y(_05217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11254_ (.Y(_05218_),
    .A(_05217_),
    .B(net1635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11255_ (.Y(_05219_),
    .B1(\acc_sum.exp_mant_logic0.a[0] ),
    .B2(net1680),
    .A2(\acc_sum.op_sign_logic0.mantisa_a[3] ),
    .A1(net1759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11256_ (.Y(_01087_),
    .A(_05218_),
    .B(_05219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11257_ (.Y(_05220_),
    .A(net1661),
    .B(\acc_sum.exp_mant_logic0.a[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11258_ (.B1(_05220_),
    .VDD(VPWR),
    .Y(_05221_),
    .VSS(VGND),
    .A1(_02959_),
    .A2(_05143_));
 sg13g2_inv_1 _11259_ (.VDD(VPWR),
    .Y(_05222_),
    .A(_05124_),
    .VSS(VGND));
 sg13g2_nand2_1 _11260_ (.Y(_05223_),
    .A(net1655),
    .B(\acc_sum.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11261_ (.B1(_05223_),
    .VDD(VPWR),
    .Y(_05224_),
    .VSS(VGND),
    .A1(_02963_),
    .A2(_05222_));
 sg13g2_nor2_1 _11262_ (.A(_05221_),
    .B(_05224_),
    .Y(_05225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11263_ (.B(_05116_),
    .C(_05020_),
    .A(_05119_),
    .Y(_05226_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05023_));
 sg13g2_nor2_2 _11264_ (.A(_05226_),
    .B(_05106_),
    .Y(_05227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11265_ (.Y(_05228_),
    .B1(_05073_),
    .B2(_05227_),
    .A2(net1808),
    .A1(_05211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11266_ (.Y(_05229_),
    .B1(net1809),
    .B2(_05192_),
    .A2(net1810),
    .A1(net1653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11267_ (.B(_05228_),
    .C(_05229_),
    .A(_05225_),
    .Y(_05230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11268_ (.Y(_05231_),
    .A(_05230_),
    .B(net1635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11269_ (.Y(_05232_),
    .A(net1761),
    .B(\acc_sum.op_sign_logic0.mantisa_a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11270_ (.Y(_01086_),
    .A(_05231_),
    .B(_05232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11271_ (.Y(_05233_),
    .A(net1655),
    .B(\acc_sum.exp_mant_logic0.a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11272_ (.Y(_05234_),
    .A(net1661),
    .B(\acc_sum.exp_mant_logic0.a[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11273_ (.Y(_05235_),
    .A(_05141_),
    .B(\acc_sum.exp_mant_logic0.a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11274_ (.B(_05234_),
    .C(_05235_),
    .A(_05233_),
    .Y(_05236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11275_ (.Y(_05237_),
    .B1(net1808),
    .B2(_05227_),
    .A2(net1809),
    .A1(_05211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11276_ (.Y(_05238_),
    .B1(net1810),
    .B2(_05192_),
    .A2(\acc_sum.exp_mant_logic0.a[3] ),
    .A1(net1653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11277_ (.Y(_05239_),
    .A(_05237_),
    .B(_05238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11278_ (.B1(net1635),
    .VDD(VPWR),
    .Y(_05240_),
    .VSS(VGND),
    .A1(_05236_),
    .A2(_05239_));
 sg13g2_nand2_1 _11279_ (.Y(_05241_),
    .A(net1761),
    .B(\acc_sum.op_sign_logic0.mantisa_a[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11280_ (.Y(_01085_),
    .A(_05240_),
    .B(_05241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11281_ (.Y(_05242_),
    .B1(net1809),
    .B2(_05227_),
    .A2(net1810),
    .A1(_05211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11282_ (.Y(_05243_),
    .B1(\acc_sum.exp_mant_logic0.a[3] ),
    .B2(_05192_),
    .A2(\acc_sum.exp_mant_logic0.a[2] ),
    .A1(net1653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11283_ (.Y(_05244_),
    .B1(\acc_sum.exp_mant_logic0.a[1] ),
    .B2(net1661),
    .A2(\acc_sum.exp_mant_logic0.a[0] ),
    .A1(_05141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11284_ (.B(_05243_),
    .C(_05244_),
    .A(_05242_),
    .Y(_05245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11285_ (.Y(_05246_),
    .A(net1635),
    .B(_05245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11286_ (.Y(_05247_),
    .A(net1761),
    .B(\acc_sum.op_sign_logic0.mantisa_a[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11287_ (.Y(_01084_),
    .A(_05246_),
    .B(_05247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11288_ (.B(_03349_),
    .C(_03355_),
    .A(_03347_),
    .Y(_05248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11289_ (.B(_03339_),
    .C(_03341_),
    .A(_03337_),
    .Y(_05249_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03343_));
 sg13g2_nand4_1 _11290_ (.B(_03331_),
    .C(_03333_),
    .A(_03329_),
    .Y(_05250_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03335_));
 sg13g2_nand4_1 _11291_ (.B(_03351_),
    .C(_03353_),
    .A(_03345_),
    .Y(_05251_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_03357_));
 sg13g2_nor4_2 _11292_ (.A(_05248_),
    .B(_05249_),
    .C(_05250_),
    .Y(_05252_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_05251_));
 sg13g2_inv_4 _11293_ (.A(_05252_),
    .Y(_05253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11294_ (.B(\acc_sum.reg1en.q[0] ),
    .C(_05253_),
    .A(_05046_),
    .Y(_05254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11295_ (.B1(_05254_),
    .VDD(VPWR),
    .Y(_01083_),
    .VSS(VGND),
    .A1(net1813),
    .A2(_02797_));
 sg13g2_a22oi_1 _11296_ (.Y(_05255_),
    .B1(_05253_),
    .B2(_05124_),
    .A2(net1697),
    .A1(net1811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _11297_ (.A(_05150_),
    .B_N(_05052_),
    .Y(_05256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_102_clk (.A(clknet_5_15__leaf_clk),
    .X(clknet_leaf_102_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11299_ (.Y(_05258_),
    .B(net1634),
    .A_N(_05255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11300_ (.Y(_05259_),
    .B1(net1811),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[9] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11301_ (.Y(_01082_),
    .A(_05258_),
    .B(_05259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11302_ (.Y(_05260_),
    .A(net1656),
    .B(_05253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11303_ (.Y(_05261_),
    .A(_05124_),
    .B(net1811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11304_ (.Y(_05262_),
    .A(net1697),
    .B(net1812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11305_ (.B(_05261_),
    .C(_05262_),
    .A(_05260_),
    .Y(_05263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11306_ (.Y(_05264_),
    .A(net1634),
    .B(_05263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11307_ (.Y(_05265_),
    .B1(net1812),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[8] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11308_ (.Y(_01081_),
    .A(_05264_),
    .B(_05265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11309_ (.Y(_05266_),
    .B1(net1812),
    .B2(_05161_),
    .A2(_05253_),
    .A1(net1654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11310_ (.Y(_05267_),
    .B1(net1811),
    .B2(net1656),
    .A2(net1697),
    .A1(\acc_sum.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11311_ (.Y(_05268_),
    .A(_05266_),
    .B(_05267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11312_ (.Y(_05269_),
    .A(net1634),
    .B(_05268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11313_ (.Y(_05270_),
    .B1(\acc_sum.exp_mant_logic0.b[4] ),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[7] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11314_ (.Y(_01080_),
    .A(_05269_),
    .B(_05270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11315_ (.Y(_05271_),
    .B1(_05146_),
    .B2(_05253_),
    .A2(net1811),
    .A1(net1654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11316_ (.Y(_05272_),
    .B1(net1812),
    .B2(net1656),
    .A2(\acc_sum.exp_mant_logic0.b[4] ),
    .A1(_05124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11317_ (.Y(_05273_),
    .A(net1697),
    .B(\acc_sum.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11318_ (.B(_05272_),
    .C(_05273_),
    .A(_05271_),
    .Y(_05274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11319_ (.Y(_05275_),
    .A(_05256_),
    .B(_05274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11320_ (.Y(_05276_),
    .B1(\acc_sum.exp_mant_logic0.b[3] ),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[6] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11321_ (.Y(_01079_),
    .A(_05275_),
    .B(_05276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11322_ (.A(_03347_),
    .B(_05143_),
    .Y(_05277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11323_ (.A(_03353_),
    .B(_05026_),
    .Y(_05278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11324_ (.A(_03351_),
    .B(_05176_),
    .Y(_05279_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11325_ (.A(_05277_),
    .B(_05278_),
    .C(_05279_),
    .Y(_05280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11326_ (.A(_05252_),
    .B(_05183_),
    .Y(_05281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11327_ (.A(_03349_),
    .B(_05173_),
    .Y(_05282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11328_ (.A(_03345_),
    .B(_05148_),
    .Y(_05283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11329_ (.A(_05281_),
    .B(_05282_),
    .C(_05283_),
    .Y(_05284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11330_ (.Y(_05285_),
    .A(_05280_),
    .B(_05284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11331_ (.Y(_05286_),
    .A(net1634),
    .B(_05285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11332_ (.Y(_05287_),
    .B1(\acc_sum.exp_mant_logic0.b[2] ),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[5] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11333_ (.Y(_01078_),
    .A(_05286_),
    .B(_05287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11334_ (.A(_03347_),
    .B(_05148_),
    .Y(_05288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11335_ (.A(_05252_),
    .B(_05194_),
    .Y(_05289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11336_ (.A(_03351_),
    .B(_05173_),
    .Y(_05290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11337_ (.A(_05288_),
    .B(_05289_),
    .C(_05290_),
    .Y(_05291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11338_ (.Y(_05292_),
    .B1(\acc_sum.exp_mant_logic0.b[2] ),
    .B2(_05161_),
    .A2(net1697),
    .A1(\acc_sum.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11339_ (.Y(_05293_),
    .B1(net1811),
    .B2(net1653),
    .A2(\acc_sum.exp_mant_logic0.b[4] ),
    .A1(net1654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11340_ (.B(_05292_),
    .C(_05293_),
    .A(_05291_),
    .Y(_05294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11341_ (.Y(_05295_),
    .A(_05294_),
    .B(net1634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11342_ (.Y(_05296_),
    .B1(\acc_sum.exp_mant_logic0.b[1] ),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[4] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11343_ (.Y(_01077_),
    .A(_05295_),
    .B(_05296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11344_ (.Y(_05297_),
    .A(net1654),
    .B(\acc_sum.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11345_ (.Y(_05298_),
    .A(net1656),
    .B(\acc_sum.exp_mant_logic0.b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11346_ (.Y(_05299_),
    .A(net1697),
    .B(\acc_sum.exp_mant_logic0.b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _11347_ (.X(_05300_),
    .A(_05297_),
    .B(_05298_),
    .C(_05299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11348_ (.Y(_05301_),
    .A(_05211_),
    .B(_05253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11349_ (.Y(_05302_),
    .A(_05181_),
    .B(net1812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11350_ (.Y(_05303_),
    .A(_05301_),
    .B(_05302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11351_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1811),
    .A2(_05192_),
    .Y(_05304_),
    .B1(_05303_));
 sg13g2_a22oi_1 _11352_ (.Y(_05305_),
    .B1(\acc_sum.exp_mant_logic0.b[1] ),
    .B2(_05161_),
    .A2(_05146_),
    .A1(\acc_sum.exp_mant_logic0.b[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11353_ (.B(_05304_),
    .C(_05305_),
    .A(_05300_),
    .Y(_05306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11354_ (.Y(_05307_),
    .A(_05306_),
    .B(net1634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11355_ (.Y(_05308_),
    .B1(\acc_sum.exp_mant_logic0.b[0] ),
    .B2(net1681),
    .A2(\acc_sum.op_sign_logic0.mantisa_b[3] ),
    .A1(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11356_ (.Y(_01076_),
    .A(_05307_),
    .B(_05308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11357_ (.Y(_05309_),
    .A(net1656),
    .B(\acc_sum.exp_mant_logic0.b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11358_ (.B1(_05309_),
    .VDD(VPWR),
    .Y(_05310_),
    .VSS(VGND),
    .A1(_03357_),
    .A2(_05222_));
 sg13g2_nand2_1 _11359_ (.Y(_05311_),
    .A(_05146_),
    .B(\acc_sum.exp_mant_logic0.b[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11360_ (.B1(_05311_),
    .VDD(VPWR),
    .Y(_05312_),
    .VSS(VGND),
    .A1(_03353_),
    .A2(_05143_));
 sg13g2_nor2_1 _11361_ (.A(_05310_),
    .B(_05312_),
    .Y(_05313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11362_ (.Y(_05314_),
    .B1(_05227_),
    .B2(_05253_),
    .A2(net1811),
    .A1(_05211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11363_ (.Y(_05315_),
    .B1(net1812),
    .B2(_05192_),
    .A2(\acc_sum.exp_mant_logic0.b[4] ),
    .A1(_05181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11364_ (.B(_05314_),
    .C(_05315_),
    .A(_05313_),
    .Y(_05316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11365_ (.Y(_05317_),
    .A(_05316_),
    .B(_05256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11366_ (.Y(_05318_),
    .A(net1761),
    .B(\acc_sum.op_sign_logic0.mantisa_b[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11367_ (.Y(_01075_),
    .A(_05317_),
    .B(_05318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11368_ (.Y(_05319_),
    .A(_05211_),
    .B(net1812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11369_ (.B1(_05319_),
    .VDD(VPWR),
    .Y(_05320_),
    .VSS(VGND),
    .A1(_03351_),
    .A2(_05183_));
 sg13g2_nor2_1 _11370_ (.A(_03349_),
    .B(_05194_),
    .Y(_05321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11371_ (.A(_03357_),
    .B(_05173_),
    .Y(_05322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11372_ (.A(_03353_),
    .B(_05148_),
    .Y(_05323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11373_ (.A(_05321_),
    .B(_05322_),
    .C(_05323_),
    .Y(_05324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11374_ (.A(_03355_),
    .B(_05143_),
    .Y(_05325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11375_ (.Y(_05326_),
    .A(_05227_),
    .B(\acc_sum.exp_mant_logic0.b[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _11376_ (.A(_05325_),
    .B_N(_05326_),
    .Y(_05327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _11377_ (.B(_05324_),
    .C(_05327_),
    .Y(_05328_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05320_));
 sg13g2_nand2_1 _11378_ (.Y(_05329_),
    .A(_05328_),
    .B(net1634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11379_ (.Y(_05330_),
    .A(net1762),
    .B(\acc_sum.op_sign_logic0.mantisa_b[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11380_ (.Y(_01074_),
    .A(_05329_),
    .B(_05330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11381_ (.Y(_05331_),
    .B1(net1812),
    .B2(_05227_),
    .A2(\acc_sum.exp_mant_logic0.b[4] ),
    .A1(_05211_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11382_ (.Y(_05332_),
    .B1(\acc_sum.exp_mant_logic0.b[3] ),
    .B2(_05192_),
    .A2(\acc_sum.exp_mant_logic0.b[2] ),
    .A1(_05181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11383_ (.Y(_05333_),
    .B1(\acc_sum.exp_mant_logic0.b[1] ),
    .B2(_05146_),
    .A2(\acc_sum.exp_mant_logic0.b[0] ),
    .A1(net1654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11384_ (.B(_05332_),
    .C(_05333_),
    .A(_05331_),
    .Y(_05334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11385_ (.Y(_05335_),
    .A(_05256_),
    .B(_05334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11386_ (.Y(_05336_),
    .A(net1761),
    .B(\acc_sum.op_sign_logic0.mantisa_b[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11387_ (.Y(_01073_),
    .A(_05335_),
    .B(_05336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11388_ (.VDD(VPWR),
    .Y(_05337_),
    .A(\fpdiv.div_out[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11389_ (.Y(_05338_),
    .A(net1707),
    .B(\fpdiv.div_out[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11390_ (.B1(_05338_),
    .VDD(VPWR),
    .Y(_01072_),
    .VSS(VGND),
    .A1(_05337_),
    .A2(net1706));
 sg13g2_inv_2 _11391_ (.Y(_05339_),
    .A(\fpdiv.div_out[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11392_ (.Y(_05340_),
    .A(net1707),
    .B(\fpdiv.div_out[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11393_ (.B1(_05340_),
    .VDD(VPWR),
    .Y(_01071_),
    .VSS(VGND),
    .A1(_05339_),
    .A2(net1706));
 sg13g2_nand2_1 _11394_ (.Y(_05341_),
    .A(net1718),
    .B(\fpdiv.div_out[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11395_ (.B1(_05341_),
    .VDD(VPWR),
    .Y(_01070_),
    .VSS(VGND),
    .A1(_05339_),
    .A2(\fpdiv.divider0.en_r ));
 sg13g2_inv_2 _11396_ (.Y(_05342_),
    .A(\fpdiv.div_out[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11397_ (.Y(_05343_),
    .A(net1707),
    .B(\fpdiv.div_out[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11398_ (.B1(_05343_),
    .VDD(VPWR),
    .Y(_01069_),
    .VSS(VGND),
    .A1(_05342_),
    .A2(net1706));
 sg13g2_nand2_1 _11399_ (.Y(_05344_),
    .A(net1718),
    .B(\fpdiv.div_out[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11400_ (.B1(_05344_),
    .VDD(VPWR),
    .Y(_01068_),
    .VSS(VGND),
    .A1(_05342_),
    .A2(\fpdiv.divider0.en_r ));
 sg13g2_inv_1 _11401_ (.VDD(VPWR),
    .Y(_05345_),
    .A(\fpdiv.div_out[5] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11402_ (.Y(_05346_),
    .A(net1707),
    .B(\fpdiv.div_out[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11403_ (.B1(_05346_),
    .VDD(VPWR),
    .Y(_01067_),
    .VSS(VGND),
    .A1(_05345_),
    .A2(net1706));
 sg13g2_nand2_1 _11404_ (.Y(_05347_),
    .A(net1718),
    .B(\fpdiv.div_out[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11405_ (.B1(_05347_),
    .VDD(VPWR),
    .Y(_01066_),
    .VSS(VGND),
    .A1(_05345_),
    .A2(\fpdiv.divider0.en_r ));
 sg13g2_inv_1 _11406_ (.VDD(VPWR),
    .Y(_05348_),
    .A(\fpdiv.div_out[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11407_ (.Y(_05349_),
    .A(net1707),
    .B(\fpdiv.div_out[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11408_ (.B1(_05349_),
    .VDD(VPWR),
    .Y(_01065_),
    .VSS(VGND),
    .A1(_05348_),
    .A2(net1706));
 sg13g2_inv_1 _11409_ (.VDD(VPWR),
    .Y(_05350_),
    .A(\fpdiv.div_out[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11410_ (.Y(_05351_),
    .A(net1707),
    .B(\fpdiv.div_out[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11411_ (.B1(_05351_),
    .VDD(VPWR),
    .Y(_01064_),
    .VSS(VGND),
    .A1(_05350_),
    .A2(net1706));
 sg13g2_nand2_1 _11412_ (.Y(_05352_),
    .A(net1718),
    .B(\fpdiv.div_out[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11413_ (.B1(_05352_),
    .VDD(VPWR),
    .Y(_01063_),
    .VSS(VGND),
    .A1(_05350_),
    .A2(\fpdiv.divider0.en_r ));
 sg13g2_inv_1 _11414_ (.VDD(VPWR),
    .Y(_05353_),
    .A(\fpdiv.div_out[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11415_ (.Y(_05354_),
    .A(net1707),
    .B(\fpdiv.div_out[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11416_ (.B1(_05354_),
    .VDD(VPWR),
    .Y(_01062_),
    .VSS(VGND),
    .A1(_05353_),
    .A2(net1706));
 sg13g2_nand2_1 _11417_ (.Y(_05355_),
    .A(net1647),
    .B(net1718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11418_ (.B1(_05355_),
    .VDD(VPWR),
    .Y(_01061_),
    .VSS(VGND),
    .A1(_05353_),
    .A2(\fpdiv.divider0.en_r ));
 sg13g2_nor2_1 _11419_ (.A(\fpdiv.reg_a_out[15] ),
    .B(net1942),
    .Y(_05356_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11420_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03327_),
    .A2(net1942),
    .Y(_01060_),
    .B1(_05356_));
 sg13g2_inv_2 _11421_ (.Y(_05357_),
    .A(\acc_sub.x2[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11422_ (.A(net1939),
    .B(\fpdiv.reg_a_out[14] ),
    .Y(_05358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11423_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05357_),
    .A2(net1939),
    .Y(_01059_),
    .B1(_05358_));
 sg13g2_inv_2 _11424_ (.Y(_05359_),
    .A(\acc_sub.x2[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11425_ (.A(net1940),
    .B(\fpdiv.reg_a_out[13] ),
    .Y(_05360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11426_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05359_),
    .A2(net1940),
    .Y(_01058_),
    .B1(_05360_));
 sg13g2_inv_1 _11427_ (.VDD(VPWR),
    .Y(_05361_),
    .A(\fpdiv.reg_a_out[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11428_ (.Y(_05362_),
    .A(\acc_sub.x2[12] ),
    .B(net1938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11429_ (.B1(_05362_),
    .VDD(VPWR),
    .Y(_01057_),
    .VSS(VGND),
    .A1(net1938),
    .A2(_05361_));
 sg13g2_inv_1 _11430_ (.VDD(VPWR),
    .Y(_05363_),
    .A(\fpdiv.reg_a_out[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11431_ (.Y(_05364_),
    .A(\acc_sub.x2[11] ),
    .B(net1938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11432_ (.B1(_05364_),
    .VDD(VPWR),
    .Y(_01056_),
    .VSS(VGND),
    .A1(net1938),
    .A2(_05363_));
 sg13g2_inv_1 _11433_ (.VDD(VPWR),
    .Y(_05365_),
    .A(\fpdiv.reg_a_out[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11434_ (.Y(_05366_),
    .A(\acc_sub.x2[10] ),
    .B(net1937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11435_ (.B1(_05366_),
    .VDD(VPWR),
    .Y(_01055_),
    .VSS(VGND),
    .A1(net1937),
    .A2(_05365_));
 sg13g2_inv_2 _11436_ (.Y(_05367_),
    .A(\acc_sub.x2[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11437_ (.A(net1937),
    .B(\fpdiv.reg_a_out[9] ),
    .Y(_05368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11438_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05367_),
    .A2(net1937),
    .Y(_01054_),
    .B1(_05368_));
 sg13g2_nor2_1 _11439_ (.A(net1940),
    .B(\fpdiv.reg_a_out[8] ),
    .Y(_05369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11440_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03601_),
    .A2(net1940),
    .Y(_01053_),
    .B1(_05369_));
 sg13g2_inv_1 _11441_ (.VDD(VPWR),
    .Y(_05370_),
    .A(\fpdiv.reg_a_out[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11442_ (.Y(_05371_),
    .A(\acc_sub.x2[7] ),
    .B(\fpdiv.reg1en.d[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11443_ (.B1(_05371_),
    .VDD(VPWR),
    .Y(_01052_),
    .VSS(VGND),
    .A1(net1944),
    .A2(_05370_));
 sg13g2_inv_1 _11444_ (.VDD(VPWR),
    .Y(_05372_),
    .A(\fpdiv.divider0.dividend[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11445_ (.Y(_05373_),
    .A(\acc_sub.x2[6] ),
    .B(net1946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11446_ (.B1(_05373_),
    .VDD(VPWR),
    .Y(_01051_),
    .VSS(VGND),
    .A1(net1947),
    .A2(_05372_));
 sg13g2_inv_1 _11447_ (.VDD(VPWR),
    .Y(_05374_),
    .A(\fpdiv.divider0.dividend[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11448_ (.Y(_05375_),
    .A(\acc_sub.x2[5] ),
    .B(net1946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11449_ (.B1(_05375_),
    .VDD(VPWR),
    .Y(_01050_),
    .VSS(VGND),
    .A1(net1947),
    .A2(_05374_));
 sg13g2_inv_1 _11450_ (.VDD(VPWR),
    .Y(_05376_),
    .A(\fpdiv.divider0.dividend[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11451_ (.Y(_05377_),
    .A(\acc_sub.x2[4] ),
    .B(net1946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11452_ (.B1(_05377_),
    .VDD(VPWR),
    .Y(_01049_),
    .VSS(VGND),
    .A1(net1946),
    .A2(_05376_));
 sg13g2_inv_1 _11453_ (.VDD(VPWR),
    .Y(_05378_),
    .A(\fpdiv.divider0.dividend[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11454_ (.Y(_05379_),
    .A(\acc_sub.x2[3] ),
    .B(net1947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11455_ (.B1(_05379_),
    .VDD(VPWR),
    .Y(_01048_),
    .VSS(VGND),
    .A1(net1947),
    .A2(_05378_));
 sg13g2_inv_1 _11456_ (.VDD(VPWR),
    .Y(_05380_),
    .A(\fpdiv.divider0.dividend[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11457_ (.Y(_05381_),
    .A(\acc_sub.x2[2] ),
    .B(net1946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11458_ (.B1(_05381_),
    .VDD(VPWR),
    .Y(_01047_),
    .VSS(VGND),
    .A1(net1947),
    .A2(_05380_));
 sg13g2_inv_2 _11459_ (.Y(_05382_),
    .A(\acc_sub.x2[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11460_ (.A(net1946),
    .B(\fpdiv.divider0.dividend[5] ),
    .Y(_05383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11461_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05382_),
    .A2(net1944),
    .Y(_01046_),
    .B1(_05383_));
 sg13g2_nand2_1 _11462_ (.Y(_05384_),
    .A(\acc_sub.x2[0] ),
    .B(net1947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11463_ (.B1(_05384_),
    .VDD(VPWR),
    .Y(_01045_),
    .VSS(VGND),
    .A1(net1947),
    .A2(_02722_));
 sg13g2_mux2_1 _11464_ (.A0(\fpdiv.reg_b_out[15] ),
    .A1(\fp16_res_pipe.x2[15] ),
    .S(net1942),
    .X(_01044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11465_ (.A0(\fpdiv.reg_b_out[14] ),
    .A1(\fp16_res_pipe.x2[14] ),
    .S(net1942),
    .X(_01043_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11466_ (.VDD(VPWR),
    .Y(_05385_),
    .A(\fpdiv.reg_b_out[13] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11467_ (.Y(_05386_),
    .A(\fp16_res_pipe.x2[13] ),
    .B(net1939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11468_ (.B1(_05386_),
    .VDD(VPWR),
    .Y(_01042_),
    .VSS(VGND),
    .A1(net1942),
    .A2(_05385_));
 sg13g2_mux2_1 _11469_ (.A0(\fpdiv.reg_b_out[12] ),
    .A1(\fp16_res_pipe.x2[12] ),
    .S(net1939),
    .X(_01041_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11470_ (.A0(\fpdiv.reg_b_out[11] ),
    .A1(\fp16_res_pipe.x2[11] ),
    .S(net1940),
    .X(_01040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11471_ (.A0(\fpdiv.reg_b_out[10] ),
    .A1(\fp16_res_pipe.x2[10] ),
    .S(net1940),
    .X(_01039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11472_ (.VDD(VPWR),
    .Y(_05387_),
    .A(\fpdiv.reg_b_out[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11473_ (.Y(_05388_),
    .A(\fp16_res_pipe.x2[9] ),
    .B(net1940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11474_ (.B1(_05388_),
    .VDD(VPWR),
    .Y(_01038_),
    .VSS(VGND),
    .A1(net1937),
    .A2(_05387_));
 sg13g2_inv_1 _11475_ (.VDD(VPWR),
    .Y(_05389_),
    .A(\fpdiv.reg_b_out[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11476_ (.Y(_05390_),
    .A(\fp16_res_pipe.x2[8] ),
    .B(net1942),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11477_ (.B1(_05390_),
    .VDD(VPWR),
    .Y(_01037_),
    .VSS(VGND),
    .A1(net1937),
    .A2(_05389_));
 sg13g2_inv_1 _11478_ (.VDD(VPWR),
    .Y(_05391_),
    .A(\fpdiv.reg_b_out[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11479_ (.Y(_05392_),
    .A(\fp16_res_pipe.x2[7] ),
    .B(\fpdiv.reg1en.d[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11480_ (.B1(_05392_),
    .VDD(VPWR),
    .Y(_01036_),
    .VSS(VGND),
    .A1(\fpdiv.reg1en.d[0] ),
    .A2(_05391_));
 sg13g2_inv_1 _11481_ (.VDD(VPWR),
    .Y(_05393_),
    .A(\fpdiv.divider0.divisor[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11482_ (.Y(_05394_),
    .A(\fp16_res_pipe.x2[6] ),
    .B(net1948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11483_ (.B1(_05394_),
    .VDD(VPWR),
    .Y(_01035_),
    .VSS(VGND),
    .A1(net1948),
    .A2(_05393_));
 sg13g2_nand2_1 _11484_ (.Y(_05395_),
    .A(\fp16_res_pipe.x2[5] ),
    .B(net1945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11485_ (.B1(_05395_),
    .VDD(VPWR),
    .Y(_01034_),
    .VSS(VGND),
    .A1(net1945),
    .A2(_01763_));
 sg13g2_nand2_1 _11486_ (.Y(_05396_),
    .A(\fp16_res_pipe.x2[4] ),
    .B(net1945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11487_ (.B1(_05396_),
    .VDD(VPWR),
    .Y(_01033_),
    .VSS(VGND),
    .A1(net1945),
    .A2(_01766_));
 sg13g2_nand2_1 _11488_ (.Y(_05397_),
    .A(\fp16_res_pipe.x2[3] ),
    .B(net1945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11489_ (.B1(_05397_),
    .VDD(VPWR),
    .Y(_01032_),
    .VSS(VGND),
    .A1(net1945),
    .A2(_01768_));
 sg13g2_mux2_1 _11490_ (.A0(\fpdiv.divider0.divisor[6] ),
    .A1(\fp16_res_pipe.x2[2] ),
    .S(net1945),
    .X(_01031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11491_ (.A0(\fpdiv.divider0.divisor[5] ),
    .A1(\fp16_res_pipe.x2[1] ),
    .S(net1944),
    .X(_01030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11492_ (.A0(\fpdiv.divider0.divisor[4] ),
    .A1(\fp16_res_pipe.x2[0] ),
    .S(net1944),
    .X(_01029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11493_ (.VDD(VPWR),
    .Y(_05398_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11494_ (.Y(_05399_),
    .A(net1840),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11495_ (.B1(_05399_),
    .VDD(VPWR),
    .Y(_05400_),
    .VSS(VGND),
    .A1(net1841),
    .A2(_05398_));
 sg13g2_inv_1 _11496_ (.VDD(VPWR),
    .Y(_05401_),
    .A(_05400_),
    .VSS(VGND));
 sg13g2_inv_1 _11497_ (.VDD(VPWR),
    .Y(_05402_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[5] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11498_ (.Y(_05403_),
    .A(net1841),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11499_ (.B1(_05403_),
    .VDD(VPWR),
    .Y(_05404_),
    .VSS(VGND),
    .A1(net1841),
    .A2(_05402_));
 sg13g2_inv_1 _11500_ (.VDD(VPWR),
    .Y(_05405_),
    .A(_05404_),
    .VSS(VGND));
 sg13g2_nand2_1 _11501_ (.Y(_05406_),
    .A(net1840),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11502_ (.VDD(VPWR),
    .Y(_05407_),
    .A(_05406_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11503_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04465_),
    .A2(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .Y(_05408_),
    .B1(_05407_));
 sg13g2_inv_2 _11504_ (.Y(_05409_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11505_ (.Y(_05410_),
    .A(net1840),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11506_ (.B1(_05410_),
    .VDD(VPWR),
    .Y(_05411_),
    .VSS(VGND),
    .A1(net1840),
    .A2(_05409_));
 sg13g2_inv_2 _11507_ (.Y(_05412_),
    .A(_05411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11508_ (.Y(_05413_),
    .A(net1840),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11509_ (.VDD(VPWR),
    .Y(_05414_),
    .A(_05413_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11510_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04465_),
    .A2(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .Y(_05415_),
    .B1(_05414_));
 sg13g2_nor2_1 _11511_ (.A(_05412_),
    .B(_05415_),
    .Y(_05416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _11512_ (.Y(_05417_),
    .B(_05416_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05408_));
 sg13g2_nor2_1 _11513_ (.A(_05405_),
    .B(_05417_),
    .Y(_05418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11514_ (.Y(_05419_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11515_ (.Y(_05420_),
    .A(net1841),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11516_ (.B1(_05420_),
    .VDD(VPWR),
    .Y(_05421_),
    .VSS(VGND),
    .A1(net1841),
    .A2(_05419_));
 sg13g2_buf_2 fanout70 (.A(net71),
    .X(net70),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11518_ (.Y(_05423_),
    .A(_05418_),
    .B(_05421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11519_ (.Y(_05424_),
    .A(_05401_),
    .B(_05423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11520_ (.VDD(VPWR),
    .Y(_05425_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .VSS(VGND));
 sg13g2_nand2_2 _11521_ (.Y(_05426_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _11522_ (.A(_05402_),
    .B(_05425_),
    .C(_05426_),
    .Y(_05427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11523_ (.Y(_05428_),
    .A(_05419_),
    .B(_05427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout86 (.A(net93),
    .X(net86),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11525_ (.VDD(VPWR),
    .Y(_05430_),
    .A(_05428_),
    .VSS(VGND));
 sg13g2_o21ai_1 _11526_ (.B1(\fp16_sum_pipe.add_renorm0.mantisa[2] ),
    .VDD(VPWR),
    .Y(_05431_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.add_renorm0.mantisa[1] ),
    .A2(\fp16_sum_pipe.add_renorm0.mantisa[0] ));
 sg13g2_inv_1 _11527_ (.VDD(VPWR),
    .Y(_05432_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _11528_ (.VDD(VPWR),
    .Y(_05433_),
    .A(_05426_),
    .VSS(VGND));
 sg13g2_a21oi_2 _11529_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_05433_),
    .Y(_05434_),
    .A2(_05432_),
    .A1(_05431_));
 sg13g2_inv_1 _11530_ (.VDD(VPWR),
    .Y(_05435_),
    .A(_05434_),
    .VSS(VGND));
 sg13g2_inv_1 _11531_ (.VDD(VPWR),
    .Y(_05436_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[8] ),
    .VSS(VGND));
 sg13g2_nand3_1 _11532_ (.B(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .C(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[5] ),
    .Y(_05437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _11533_ (.A(_05436_),
    .B(_05398_),
    .C(_05419_),
    .D(_05437_),
    .Y(_05438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11534_ (.Y(_05439_),
    .A(_05431_),
    .B(_05426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11535_ (.B(\fp16_sum_pipe.add_renorm0.mantisa[9] ),
    .C(_05439_),
    .A(_05438_),
    .Y(_05440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11536_ (.VDD(VPWR),
    .Y(_05441_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[10] ),
    .VSS(VGND));
 sg13g2_nand2_2 _11537_ (.Y(_05442_),
    .A(_05440_),
    .B(_05441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout96 (.A(net107),
    .X(net96),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _11539_ (.A(_05442_),
    .Y(_05444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11540_ (.Y(_05445_),
    .A(_05438_),
    .B(_05439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11541_ (.B(\fp16_sum_pipe.add_renorm0.mantisa[7] ),
    .C(\fp16_sum_pipe.add_renorm0.mantisa[6] ),
    .A(_05427_),
    .Y(_05446_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11542_ (.Y(_05447_),
    .A(_05446_),
    .B(_05436_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _11543_ (.A(_05445_),
    .B(_05447_),
    .X(_05448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11544_ (.VDD(VPWR),
    .Y(_05449_),
    .A(_05448_),
    .VSS(VGND));
 sg13g2_nand2_1 _11545_ (.Y(_05450_),
    .A(_05444_),
    .B(_05449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11546_ (.VDD(VPWR),
    .Y(_05451_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[9] ),
    .VSS(VGND));
 sg13g2_o21ai_1 _11547_ (.B1(_05445_),
    .VDD(VPWR),
    .Y(_05452_),
    .VSS(VGND),
    .A1(_05451_),
    .A2(_05409_));
 sg13g2_nand2_1 _11548_ (.Y(_05453_),
    .A(_05438_),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11549_ (.Y(_05454_),
    .A(_05452_),
    .B(_05453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11550_ (.B1(_05454_),
    .VDD(VPWR),
    .Y(_05455_),
    .VSS(VGND),
    .A1(_05451_),
    .A2(_05439_));
 sg13g2_buf_2 fanout118 (.A(net119),
    .X(net118),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11552_ (.A(_05450_),
    .B(_05455_),
    .Y(_05457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _11553_ (.A2(\fp16_sum_pipe.add_renorm0.mantisa[6] ),
    .A1(_05427_),
    .B1(\fp16_sum_pipe.add_renorm0.mantisa[7] ),
    .X(_05458_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _11554_ (.A(_05458_),
    .B(_05446_),
    .X(_05459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout97 (.A(net100),
    .X(net97),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11556_ (.VDD(VPWR),
    .Y(_05461_),
    .A(_05459_),
    .VSS(VGND));
 sg13g2_nand2_2 _11557_ (.Y(_05462_),
    .A(_05457_),
    .B(_05461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11558_ (.A(_05430_),
    .B(_05435_),
    .C(_05462_),
    .Y(_05463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11559_ (.VDD(VPWR),
    .Y(_05464_),
    .A(_05455_),
    .VSS(VGND));
 sg13g2_nor2_2 _11560_ (.A(_05442_),
    .B(_05464_),
    .Y(_05465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11562_ (.Y(_05467_),
    .B1(_05428_),
    .B2(_05465_),
    .A2(_05459_),
    .A1(_05442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11563_ (.Y(_05468_),
    .A(_05457_),
    .B(_05459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11564_ (.VDD(VPWR),
    .Y(_05469_),
    .A(_05468_),
    .VSS(VGND));
 sg13g2_xnor2_1 _11565_ (.Y(_05470_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .B(_05426_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout71 (.A(net72),
    .X(net71),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11567_ (.Y(_05472_),
    .A(_05469_),
    .B(_05470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11568_ (.A(_05442_),
    .B(_05455_),
    .Y(_05473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11569_ (.Y(_05474_),
    .A(_05473_),
    .B(_05448_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11570_ (.Y(_05475_),
    .A(_05474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11571_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05433_),
    .A2(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .Y(_05476_),
    .B1(\fp16_sum_pipe.add_renorm0.mantisa[5] ));
 sg13g2_nor2_2 _11572_ (.A(_05427_),
    .B(_05476_),
    .Y(_05477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11573_ (.Y(_05478_),
    .A(_05475_),
    .B(_05477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11574_ (.B(_05472_),
    .C(_05478_),
    .A(_05467_),
    .Y(_05479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11575_ (.B1(net1836),
    .VDD(VPWR),
    .Y(_05480_),
    .VSS(VGND),
    .A1(_05463_),
    .A2(_05479_));
 sg13g2_o21ai_1 _11576_ (.B1(_05480_),
    .VDD(VPWR),
    .Y(_05481_),
    .VSS(VGND),
    .A1(net1837),
    .A2(_05424_));
 sg13g2_inv_1 _11577_ (.VDD(VPWR),
    .Y(_05482_),
    .A(_05477_),
    .VSS(VGND));
 sg13g2_nor3_2 _11578_ (.A(_05428_),
    .B(_05482_),
    .C(_05462_),
    .Y(_05483_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11579_ (.A(_05477_),
    .B(_05428_),
    .Y(_05484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11580_ (.VDD(VPWR),
    .Y(_05485_),
    .A(_05484_),
    .VSS(VGND));
 sg13g2_nor4_1 _11581_ (.A(_05485_),
    .B(_05470_),
    .C(_05435_),
    .D(_05462_),
    .Y(_05486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11582_ (.A(_05469_),
    .B(_05486_),
    .Y(_05487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11583_ (.Y(_05488_),
    .A(_05487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _11584_ (.A(_05483_),
    .B(_05465_),
    .C(_05488_),
    .Y(_05489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11585_ (.B(_05449_),
    .C(_05461_),
    .A(_05464_),
    .Y(_05490_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05428_));
 sg13g2_nand2_2 _11586_ (.Y(_05491_),
    .A(_05490_),
    .B(_05444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _11587_ (.X(_05492_),
    .A(_05461_),
    .B(_05484_),
    .C(_05470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _11588_ (.Y(_05493_),
    .A(_05457_),
    .B(_05492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11589_ (.VDD(VPWR),
    .Y(_05494_),
    .A(_05493_),
    .VSS(VGND));
 sg13g2_nor2_2 _11590_ (.A(_05475_),
    .B(_05494_),
    .Y(_05495_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _11591_ (.A(_05495_),
    .Y(_05496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11592_ (.A(_05491_),
    .B(_05496_),
    .Y(_05497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11593_ (.Y(_05498_),
    .A(net1836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1769 (.A(_03740_),
    .X(net1769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11595_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05489_),
    .A2(_05497_),
    .Y(_05500_),
    .B1(net1757));
 sg13g2_nand2_1 _11596_ (.Y(_05501_),
    .A(net1841),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11597_ (.B1(_05501_),
    .VDD(VPWR),
    .Y(_05502_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .A2(_05436_));
 sg13g2_nor2_1 _11598_ (.A(_05401_),
    .B(_05423_),
    .Y(_05503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11599_ (.B(_05421_),
    .C(_05400_),
    .A(_05418_),
    .Y(_05504_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05502_));
 sg13g2_o21ai_1 _11600_ (.B1(_05504_),
    .VDD(VPWR),
    .Y(_05505_),
    .VSS(VGND),
    .A1(_05502_),
    .A2(_05503_));
 sg13g2_nor2_1 _11601_ (.A(_05430_),
    .B(_05462_),
    .Y(_05506_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11602_ (.A(_05482_),
    .B(_05468_),
    .Y(_05507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11603_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05506_),
    .A2(_05470_),
    .Y(_05508_),
    .B1(_05507_));
 sg13g2_nand2_1 _11604_ (.Y(_05509_),
    .A(_05483_),
    .B(_05434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11605_ (.Y(_05510_),
    .A(_05465_),
    .B(_05459_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11606_ (.A(_05449_),
    .B(_05444_),
    .Y(_05511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11607_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05475_),
    .A2(_05428_),
    .Y(_05512_),
    .B1(_05511_));
 sg13g2_nand4_1 _11608_ (.B(_05509_),
    .C(_05510_),
    .A(_05508_),
    .Y(_05513_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05512_));
 sg13g2_nand2_1 _11609_ (.Y(_05514_),
    .A(_05513_),
    .B(net1836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11610_ (.B1(_05514_),
    .VDD(VPWR),
    .Y(_05515_),
    .VSS(VGND),
    .A1(net1836),
    .A2(_05505_));
 sg13g2_nor3_1 _11611_ (.A(_05481_),
    .B(_05500_),
    .C(_05515_),
    .Y(_05516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11612_ (.VDD(VPWR),
    .Y(_05517_),
    .A(_05415_),
    .VSS(VGND));
 sg13g2_nor2_1 _11613_ (.A(net1840),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[0] ),
    .Y(_05518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1840),
    .A2(_05409_),
    .Y(_05519_),
    .B1(_05518_));
 sg13g2_nor3_1 _11615_ (.A(\fp16_sum_pipe.add_renorm0.mantisa[1] ),
    .B(_05519_),
    .C(_05412_),
    .Y(_05520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11616_ (.A(_05412_),
    .B(_05520_),
    .Y(_05521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11617_ (.VDD(VPWR),
    .Y(_05522_),
    .A(_05416_),
    .VSS(VGND));
 sg13g2_o21ai_1 _11618_ (.B1(_05522_),
    .VDD(VPWR),
    .Y(_05523_),
    .VSS(VGND),
    .A1(_05517_),
    .A2(_05521_));
 sg13g2_nand2_1 _11619_ (.Y(_05524_),
    .A(_05523_),
    .B(net1757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11620_ (.A(net1838),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[10] ),
    .Y(_05525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11621_ (.VDD(VPWR),
    .Y(_05526_),
    .A(_05525_),
    .VSS(VGND));
 sg13g2_nand2_1 _11622_ (.Y(_05527_),
    .A(_05421_),
    .B(_05404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _11623_ (.A(_05401_),
    .B(_05415_),
    .C(_05408_),
    .D(_05527_),
    .Y(_05528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11624_ (.Y(_05529_),
    .A(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .B(\fp16_sum_pipe.add_renorm0.mantisa[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11625_ (.B1(_05529_),
    .VDD(VPWR),
    .Y(_05530_),
    .VSS(VGND),
    .A1(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .A2(_05451_));
 sg13g2_nand3_1 _11626_ (.B(_05502_),
    .C(_05530_),
    .A(_05528_),
    .Y(_05531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11627_ (.Y(_05532_),
    .A(_05526_),
    .B(_05531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11628_ (.Y(_05533_),
    .A(_05532_),
    .B(_05520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11629_ (.Y(_05534_),
    .A(_05532_),
    .B(_05521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11630_ (.A(_05416_),
    .B(_05521_),
    .Y(_05535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _11631_ (.A(_05535_),
    .B(_05525_),
    .C(_05531_),
    .Y(_05536_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11632_ (.VDD(VPWR),
    .Y(_05537_),
    .A(_05536_),
    .VSS(VGND));
 sg13g2_nand2_1 _11633_ (.Y(_05538_),
    .A(_05412_),
    .B(_05526_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11634_ (.B(_05534_),
    .C(_05537_),
    .A(_05533_),
    .Y(_05539_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05538_));
 sg13g2_o21ai_1 _11635_ (.B1(net1837),
    .VDD(VPWR),
    .Y(_05540_),
    .VSS(VGND),
    .A1(_05435_),
    .A2(_05444_));
 sg13g2_o21ai_1 _11636_ (.B1(_05540_),
    .VDD(VPWR),
    .Y(_05541_),
    .VSS(VGND),
    .A1(_05524_),
    .A2(_05539_));
 sg13g2_nor2_1 _11637_ (.A(_05430_),
    .B(_05468_),
    .Y(_05542_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11638_ (.Y(_05543_),
    .B1(_05470_),
    .B2(_05483_),
    .A2(_05506_),
    .A1(_05477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11639_ (.Y(_05544_),
    .B1(_05434_),
    .B2(_05494_),
    .A2(_05459_),
    .A1(_05475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11640_ (.Y(_05545_),
    .A(_05455_),
    .B(_05450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11641_ (.B(_05544_),
    .C(_05545_),
    .A(_05543_),
    .Y(_05546_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11642_ (.B1(net1836),
    .VDD(VPWR),
    .Y(_05547_),
    .VSS(VGND),
    .A1(_05542_),
    .A2(_05546_));
 sg13g2_xnor2_1 _11643_ (.Y(_05548_),
    .A(_05530_),
    .B(_05504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11644_ (.Y(_05549_),
    .A(_05548_),
    .B(_05498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11645_ (.Y(_05550_),
    .A(_05547_),
    .B(_05549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11646_ (.Y(_05551_),
    .A(_05550_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11647_ (.Y(_05552_),
    .B1(_05434_),
    .B2(_05465_),
    .A2(_05470_),
    .A1(_05442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11648_ (.Y(_05553_),
    .A(_05522_),
    .B(_05408_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11649_ (.B(_05498_),
    .C(_05417_),
    .A(_05553_),
    .Y(_05554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11650_ (.B1(_05554_),
    .VDD(VPWR),
    .Y(_05555_),
    .VSS(VGND),
    .A1(_05498_),
    .A2(_05552_));
 sg13g2_a22oi_1 _11651_ (.Y(_05556_),
    .B1(_05477_),
    .B2(_05465_),
    .A2(_05428_),
    .A1(_05442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11652_ (.Y(_05557_),
    .A(_05469_),
    .B(_05434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11653_ (.Y(_05558_),
    .A(_05475_),
    .B(_05470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11654_ (.B(_05557_),
    .C(_05558_),
    .A(_05556_),
    .Y(_05559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11655_ (.Y(_05560_),
    .A(_05421_),
    .B(_05418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11656_ (.A(net1836),
    .B(_05560_),
    .Y(_05561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11657_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05559_),
    .A2(net1837),
    .Y(_05562_),
    .B1(_05561_));
 sg13g2_inv_1 _11658_ (.VDD(VPWR),
    .Y(_05563_),
    .A(_05562_),
    .VSS(VGND));
 sg13g2_xnor2_1 _11659_ (.Y(_05564_),
    .A(_05405_),
    .B(_05417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11660_ (.Y(_05565_),
    .B1(_05470_),
    .B2(_05465_),
    .A2(_05477_),
    .A1(_05442_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11661_ (.Y(_05566_),
    .A(_05475_),
    .B(_05434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _11662_ (.A2(_05566_),
    .A1(_05565_),
    .B1(_05498_),
    .X(_05567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11663_ (.B1(_05567_),
    .VDD(VPWR),
    .Y(_05568_),
    .VSS(VGND),
    .A1(net1836),
    .A2(_05564_));
 sg13g2_nor3_1 _11664_ (.A(_05555_),
    .B(_05563_),
    .C(_05568_),
    .Y(_05569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11665_ (.B(_05541_),
    .C(_05551_),
    .A(_05516_),
    .Y(_05570_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05569_));
 sg13g2_buf_2 place1665 (.A(_01591_),
    .X(net1665),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _11667_ (.Y(_05572_),
    .A(_05570_),
    .B(\fp16_sum_pipe.reg3en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _11668_ (.A(\fp16_sum_pipe.reg3en.q[0] ),
    .Y(_05573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1774 (.A(_02179_),
    .X(net1774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11670_ (.Y(_05575_),
    .A(_05573_),
    .B(\add_result[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11671_ (.B1(_05575_),
    .VDD(VPWR),
    .Y(_01028_),
    .VSS(VGND),
    .A1(_04389_),
    .A2(_05572_));
 sg13g2_nand3_1 _11672_ (.B(\fp16_sum_pipe.add_renorm0.exp[1] ),
    .C(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .A(\fp16_sum_pipe.add_renorm0.exp[2] ),
    .Y(_05576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11673_ (.A(_04589_),
    .B(_05576_),
    .Y(_05577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11674_ (.Y(_05578_),
    .A(_05577_),
    .B(\fp16_sum_pipe.add_renorm0.exp[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11675_ (.A(_04585_),
    .B(_05578_),
    .Y(_05579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11676_ (.Y(_05580_),
    .A(_05579_),
    .B(\fp16_sum_pipe.add_renorm0.exp[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11677_ (.Y(_05581_),
    .A(_04581_),
    .B(_05580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11678_ (.VDD(VPWR),
    .Y(_05582_),
    .A(_05581_),
    .VSS(VGND));
 sg13g2_nor2_2 _11679_ (.A(_05441_),
    .B(_05440_),
    .Y(_05583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout100 (.A(net107),
    .X(net100),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout99 (.A(net100),
    .X(net99),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11682_ (.A(_04581_),
    .B(net1727),
    .Y(_05586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _11683_ (.A2(net1727),
    .A1(_05582_),
    .B1(_05586_),
    .X(_05587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1701 (.A(_06567_),
    .X(net1701),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11685_ (.Y(_05589_),
    .A(_04589_),
    .B(_05576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11686_ (.A(\fp16_sum_pipe.add_renorm0.exp[3] ),
    .B(_05583_),
    .Y(_05590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11687_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05583_),
    .A2(_05589_),
    .Y(_05591_),
    .B1(_05590_));
 sg13g2_inv_2 _11688_ (.Y(_05592_),
    .A(_05591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11689_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fp16_sum_pipe.add_renorm0.exp[1] ),
    .A2(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .Y(_05593_),
    .B1(\fp16_sum_pipe.add_renorm0.exp[2] ));
 sg13g2_nor2b_1 _11690_ (.A(_05593_),
    .B_N(_05576_),
    .Y(_05594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11691_ (.Y(_05595_),
    .A(_05583_),
    .B(_05594_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11692_ (.B1(_05595_),
    .VDD(VPWR),
    .Y(_05596_),
    .VSS(VGND),
    .A1(_04591_),
    .A2(_05583_));
 sg13g2_buf_1 fanout126 (.A(net127),
    .X(net126),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11694_ (.Y(_05598_),
    .A(_05596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11695_ (.B(_05598_),
    .C(_05444_),
    .A(_05592_),
    .Y(_05599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11697_ (.VDD(VPWR),
    .Y(_05601_),
    .A(_05599_),
    .VSS(VGND));
 sg13g2_xnor2_1 _11698_ (.Y(_05602_),
    .A(_04587_),
    .B(_05577_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11699_ (.Y(_05603_),
    .A(net1727),
    .B(_05602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11700_ (.B1(_05603_),
    .VDD(VPWR),
    .Y(_05604_),
    .VSS(VGND),
    .A1(_04587_),
    .A2(net1727));
 sg13g2_buf_1 fanout135 (.A(net136),
    .X(net135),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11702_ (.Y(_05606_),
    .A(\fp16_sum_pipe.add_renorm0.exp[5] ),
    .B(_05578_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11703_ (.Y(_05607_),
    .A(net1727),
    .B(_05606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11704_ (.B1(_05607_),
    .VDD(VPWR),
    .Y(_05608_),
    .VSS(VGND),
    .A1(_04585_),
    .A2(net1727));
 sg13g2_buf_2 fanout136 (.A(net140),
    .X(net136),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11706_ (.A(_05604_),
    .B(_05608_),
    .Y(_05610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11707_ (.Y(_05611_),
    .A(_05601_),
    .B(_05610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11708_ (.VDD(VPWR),
    .Y(_05612_),
    .A(_05611_),
    .VSS(VGND));
 sg13g2_nand2_1 _11709_ (.Y(_05613_),
    .A(_05612_),
    .B(_04583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11710_ (.Y(_05614_),
    .A(_05587_),
    .B(_05613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11711_ (.Y(_05615_),
    .A(_05583_),
    .B(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11712_ (.Y(_05616_),
    .A(\fp16_sum_pipe.add_renorm0.exp[1] ),
    .B(_05615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11713_ (.Y(_05617_),
    .A(_05616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11714_ (.Y(_05618_),
    .A(_05596_),
    .B(_05493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11715_ (.A(_05617_),
    .B(_05618_),
    .Y(_05619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05493_),
    .A2(_05596_),
    .Y(_05620_),
    .B1(_05619_));
 sg13g2_inv_2 _11717_ (.Y(_05621_),
    .A(_05604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11718_ (.B(_05621_),
    .C(_05592_),
    .A(_05620_),
    .Y(_05622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_5_21__leaf_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11720_ (.A(_05608_),
    .B(_05622_),
    .Y(_05624_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11721_ (.Y(_05625_),
    .A(\fp16_sum_pipe.add_renorm0.exp[6] ),
    .B(_05579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11722_ (.A(\fp16_sum_pipe.add_renorm0.exp[6] ),
    .B(net1727),
    .Y(_05626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _11723_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_05626_),
    .Y(_05627_),
    .A2(_05625_),
    .A1(net1727));
 sg13g2_inv_1 _11724_ (.VDD(VPWR),
    .Y(_05628_),
    .A(_05627_),
    .VSS(VGND));
 sg13g2_nand2_1 _11725_ (.Y(_05629_),
    .A(_05624_),
    .B(_05628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11726_ (.Y(_05630_),
    .A(_05587_),
    .B(_05629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _11727_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_05496_),
    .C1(net1757),
    .B1(_05630_),
    .A1(_05491_),
    .Y(_05631_),
    .A2(_05614_));
 sg13g2_nor2_1 _11728_ (.A(_05483_),
    .B(_05486_),
    .Y(_05632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11729_ (.Y(_05633_),
    .A(_05632_),
    .B(_05596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11730_ (.Y(_05634_),
    .A(_05633_),
    .B(_05592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11731_ (.Y(_05635_),
    .A(_05488_),
    .B(_05617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11732_ (.Y(_05636_),
    .A(_04595_),
    .B(_05583_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11733_ (.A(_05617_),
    .B(_05488_),
    .Y(_05637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11734_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05635_),
    .A2(_05636_),
    .Y(_05638_),
    .B1(_05637_));
 sg13g2_xnor2_1 _11735_ (.Y(_05639_),
    .A(_05596_),
    .B(_05632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11736_ (.Y(_05640_),
    .B(_05592_),
    .A_N(_05639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11737_ (.A(_05638_),
    .B(_05640_),
    .Y(_05641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _11738_ (.A(_05634_),
    .B(_05641_),
    .Y(_05642_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_52_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_52_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11740_ (.Y(_05644_),
    .A(_05642_),
    .B(_05610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11741_ (.VDD(VPWR),
    .Y(_05645_),
    .A(_05587_),
    .VSS(VGND));
 sg13g2_o21ai_1 _11742_ (.B1(_05645_),
    .VDD(VPWR),
    .Y(_05646_),
    .VSS(VGND),
    .A1(_05627_),
    .A2(_05644_));
 sg13g2_nand4_1 _11743_ (.B(_05587_),
    .C(_05628_),
    .A(_05642_),
    .Y(_05647_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05610_));
 sg13g2_inv_4 _11744_ (.A(_05489_),
    .Y(_05648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11745_ (.B(_05647_),
    .C(_05648_),
    .A(_05646_),
    .Y(_05649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11746_ (.Y(_05650_),
    .A(_05631_),
    .B(_05649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11747_ (.A(net1839),
    .B(\fp16_sum_pipe.add_renorm0.exp[7] ),
    .Y(_05651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05581_),
    .A2(net1839),
    .Y(_05652_),
    .B1(_05651_));
 sg13g2_nand2_1 _11749_ (.Y(_05653_),
    .A(_05625_),
    .B(net1839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11750_ (.B1(_05653_),
    .VDD(VPWR),
    .Y(_05654_),
    .VSS(VGND),
    .A1(net1839),
    .A2(\fp16_sum_pipe.add_renorm0.exp[6] ));
 sg13g2_nor2_1 _11751_ (.A(net1839),
    .B(_04587_),
    .Y(_05655_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11752_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05602_),
    .A2(net1839),
    .Y(_05656_),
    .B1(_05655_));
 sg13g2_nand2_1 _11753_ (.Y(_05657_),
    .A(_04465_),
    .B(\fp16_sum_pipe.add_renorm0.exp[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11754_ (.B1(_05657_),
    .VDD(VPWR),
    .Y(_05658_),
    .VSS(VGND),
    .A1(_04465_),
    .A2(_05589_));
 sg13g2_inv_1 _11755_ (.VDD(VPWR),
    .Y(_05659_),
    .A(_05658_),
    .VSS(VGND));
 sg13g2_nand2_1 _11756_ (.Y(_05660_),
    .A(_05594_),
    .B(net1838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11757_ (.B1(_05660_),
    .VDD(VPWR),
    .Y(_05661_),
    .VSS(VGND),
    .A1(net1838),
    .A2(_04591_));
 sg13g2_inv_1 _11758_ (.VDD(VPWR),
    .Y(_05662_),
    .A(_05661_),
    .VSS(VGND));
 sg13g2_nor2_1 _11759_ (.A(net1838),
    .B(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .Y(_05663_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11760_ (.Y(_05664_),
    .A(net1838),
    .B(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _11761_ (.A(_05663_),
    .B_N(_05664_),
    .Y(_05665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11762_ (.B(\fp16_sum_pipe.add_renorm0.exp[1] ),
    .C(_05665_),
    .A(_05536_),
    .Y(_05666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11763_ (.A(_05662_),
    .B(_05666_),
    .Y(_05667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11764_ (.VDD(VPWR),
    .Y(_05668_),
    .A(_05667_),
    .VSS(VGND));
 sg13g2_nor3_1 _11765_ (.A(_05656_),
    .B(_05659_),
    .C(_05668_),
    .Y(_05669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11766_ (.Y(_05670_),
    .A(_05606_),
    .B(net1839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11767_ (.B1(_05670_),
    .VDD(VPWR),
    .Y(_05671_),
    .VSS(VGND),
    .A1(net1839),
    .A2(_04585_));
 sg13g2_nand2_1 _11768_ (.Y(_05672_),
    .A(_05669_),
    .B(_05671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11769_ (.A(_05654_),
    .B(_05672_),
    .Y(_05673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11770_ (.Y(_05674_),
    .A(_05652_),
    .B(_05673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11771_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1758),
    .A2(_05674_),
    .Y(_05675_),
    .B1(_05572_));
 sg13g2_nand2_1 _11772_ (.Y(_05676_),
    .A(_05650_),
    .B(_05675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11773_ (.Y(_05677_),
    .A(_05573_),
    .B(\add_result[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11774_ (.Y(_01027_),
    .A(_05676_),
    .B(_05677_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _11775_ (.A(_05672_),
    .B(_05654_),
    .X(_05678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11776_ (.B1(net1758),
    .VDD(VPWR),
    .Y(_05679_),
    .VSS(VGND),
    .A1(_05673_),
    .A2(_05678_));
 sg13g2_nand3_1 _11777_ (.B(\fp16_sum_pipe.reg3en.q[0] ),
    .C(_05679_),
    .A(_05570_),
    .Y(_05680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11778_ (.Y(_05681_),
    .A(_05644_),
    .B(_05628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11779_ (.B(_05627_),
    .C(_05610_),
    .A(_05642_),
    .Y(_05682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11780_ (.B(_05682_),
    .C(_05648_),
    .A(_05681_),
    .Y(_05683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11781_ (.Y(_05684_),
    .A(_05611_),
    .B(_05627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11782_ (.Y(_05685_),
    .B1(_05684_),
    .B2(_05613_),
    .A2(_05490_),
    .A1(_05444_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11783_ (.VDD(VPWR),
    .Y(_05686_),
    .A(_05624_),
    .VSS(VGND));
 sg13g2_nand2_1 _11784_ (.Y(_05687_),
    .A(_05686_),
    .B(_05627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05687_),
    .A2(_05629_),
    .Y(_05688_),
    .B1(_05495_));
 sg13g2_nor3_1 _11786_ (.A(net1757),
    .B(_05685_),
    .C(_05688_),
    .Y(_05689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _11787_ (.A(_05683_),
    .B(_05689_),
    .X(_05690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11788_ (.Y(_05691_),
    .A(_05573_),
    .B(\add_result[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11789_ (.B1(_05691_),
    .VDD(VPWR),
    .Y(_01026_),
    .VSS(VGND),
    .A1(_05680_),
    .A2(_05690_));
 sg13g2_a21oi_1 _11790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05642_),
    .A2(_05621_),
    .Y(_05692_),
    .B1(_05608_));
 sg13g2_nand3_1 _11791_ (.B(_05608_),
    .C(_05621_),
    .A(_05642_),
    .Y(_05693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _11792_ (.B(_05648_),
    .C(_05693_),
    .Y(_05694_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05692_));
 sg13g2_nand2_1 _11793_ (.Y(_05695_),
    .A(_05601_),
    .B(_05621_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _11794_ (.A2(_05695_),
    .A1(_05608_),
    .B1(_05612_),
    .X(_05696_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11795_ (.Y(_05697_),
    .A(_05608_),
    .B(_05622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11796_ (.Y(_05698_),
    .B1(_05496_),
    .B2(_05697_),
    .A2(_05696_),
    .A1(_05491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11797_ (.B(net1837),
    .C(_05698_),
    .A(_05694_),
    .Y(_05699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11798_ (.Y(_05700_),
    .A(_05671_),
    .B(_05669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11799_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1758),
    .A2(_05700_),
    .Y(_05701_),
    .B1(_05572_));
 sg13g2_nand2_1 _11800_ (.Y(_05702_),
    .A(_05699_),
    .B(_05701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11801_ (.Y(_05703_),
    .A(_05573_),
    .B(\add_result[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11802_ (.Y(_01025_),
    .A(_05702_),
    .B(_05703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11803_ (.B1(_05656_),
    .VDD(VPWR),
    .Y(_05704_),
    .VSS(VGND),
    .A1(_05659_),
    .A2(_05668_));
 sg13g2_nand2b_1 _11804_ (.Y(_05705_),
    .B(_05704_),
    .A_N(_05669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11805_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1758),
    .A2(_05705_),
    .Y(_05706_),
    .B1(_05572_));
 sg13g2_o21ai_1 _11806_ (.B1(_05621_),
    .VDD(VPWR),
    .Y(_05707_),
    .VSS(VGND),
    .A1(_05634_),
    .A2(_05641_));
 sg13g2_nand2_1 _11807_ (.Y(_05708_),
    .A(_05642_),
    .B(_05604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11808_ (.B(_05708_),
    .C(_05648_),
    .A(_05707_),
    .Y(_05709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11809_ (.Y(_05710_),
    .A(_05604_),
    .B(_05599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11810_ (.Y(_05711_),
    .A(_05620_),
    .B(_05592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11811_ (.Y(_05712_),
    .A(_05711_),
    .B(_05604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11812_ (.Y(_05713_),
    .A(_05712_),
    .B(_05622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11813_ (.Y(_05714_),
    .B1(_05496_),
    .B2(_05713_),
    .A2(_05710_),
    .A1(_05491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11814_ (.B(net1837),
    .C(_05714_),
    .A(_05709_),
    .Y(_05715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11815_ (.Y(_05716_),
    .A(_05706_),
    .B(_05715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11816_ (.Y(_05717_),
    .A(_05573_),
    .B(\add_result[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11817_ (.Y(_01024_),
    .A(_05716_),
    .B(_05717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11818_ (.Y(_05718_),
    .A(_05658_),
    .B(_05667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11819_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1758),
    .A2(_05718_),
    .Y(_05719_),
    .B1(_05572_));
 sg13g2_or2_1 _11820_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_05720_),
    .B(_05638_),
    .A(_05639_));
 sg13g2_a21oi_1 _11821_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05720_),
    .A2(_05633_),
    .Y(_05721_),
    .B1(_05592_));
 sg13g2_o21ai_1 _11822_ (.B1(_05648_),
    .VDD(VPWR),
    .Y(_05722_),
    .VSS(VGND),
    .A1(_05642_),
    .A2(_05721_));
 sg13g2_a21oi_1 _11823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05598_),
    .A2(_05444_),
    .Y(_05723_),
    .B1(_05592_));
 sg13g2_nand2b_1 _11824_ (.Y(_05724_),
    .B(_05599_),
    .A_N(_05723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _11825_ (.Y(_05725_),
    .B(_05591_),
    .A_N(_05620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11826_ (.Y(_05726_),
    .A(_05725_),
    .B(_05711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _11827_ (.Y(_05727_),
    .B1(_05496_),
    .B2(_05726_),
    .A2(_05724_),
    .A1(_05491_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _11828_ (.B(net1837),
    .C(_05727_),
    .A(_05722_),
    .Y(_05728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11829_ (.Y(_05729_),
    .A(_05719_),
    .B(_05728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11830_ (.Y(_05730_),
    .A(net1756),
    .B(\add_result[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11831_ (.Y(_01023_),
    .A(_05729_),
    .B(_05730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11832_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05638_),
    .A2(_05639_),
    .Y(_05731_),
    .B1(_05489_));
 sg13g2_nand2_1 _11833_ (.Y(_05732_),
    .A(_05731_),
    .B(_05720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11834_ (.A(_05444_),
    .B(_05598_),
    .Y(_05733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11835_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05506_),
    .A2(_05598_),
    .Y(_05734_),
    .B1(_05733_));
 sg13g2_nand2_1 _11836_ (.Y(_05735_),
    .A(_05618_),
    .B(_05617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _11837_ (.B(_05496_),
    .C(_05735_),
    .Y(_05736_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05619_));
 sg13g2_nand4_1 _11838_ (.B(net1837),
    .C(_05734_),
    .A(_05732_),
    .Y(_05737_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05736_));
 sg13g2_and2_1 _11839_ (.A(_05666_),
    .B(_05662_),
    .X(_05738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11840_ (.B1(net1758),
    .VDD(VPWR),
    .Y(_05739_),
    .VSS(VGND),
    .A1(_05667_),
    .A2(_05738_));
 sg13g2_nand3_1 _11841_ (.B(_05737_),
    .C(_05739_),
    .A(_05570_),
    .Y(_05740_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11842_ (.Y(_05741_),
    .A(net1756),
    .B(\add_result[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11843_ (.B1(_05741_),
    .VDD(VPWR),
    .Y(_01022_),
    .VSS(VGND),
    .A1(net1756),
    .A2(_05740_));
 sg13g2_inv_1 _11844_ (.VDD(VPWR),
    .Y(_05742_),
    .A(_05637_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11845_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05742_),
    .A2(_05635_),
    .Y(_05743_),
    .B1(_05636_));
 sg13g2_nand3_1 _11846_ (.B(_05635_),
    .C(_05636_),
    .A(_05742_),
    .Y(_05744_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _11847_ (.B(_05648_),
    .C(_05744_),
    .Y(_05745_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05743_));
 sg13g2_nand2_1 _11848_ (.Y(_05746_),
    .A(_05491_),
    .B(_05616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11849_ (.Y(_05747_),
    .A(_05496_),
    .B(_05617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _11850_ (.B(net1837),
    .C(_05746_),
    .A(_05745_),
    .Y(_05748_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05747_));
 sg13g2_a21oi_1 _11851_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05537_),
    .A2(_05664_),
    .Y(_05749_),
    .B1(_05663_));
 sg13g2_a21oi_1 _11852_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05749_),
    .A2(_04593_),
    .Y(_05750_),
    .B1(\fp16_sum_pipe.seg_reg1.q[21] ));
 sg13g2_o21ai_1 _11853_ (.B1(_05750_),
    .VDD(VPWR),
    .Y(_05751_),
    .VSS(VGND),
    .A1(_04593_),
    .A2(_05749_));
 sg13g2_nand3_1 _11854_ (.B(_05748_),
    .C(_05751_),
    .A(_05570_),
    .Y(_05752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11855_ (.Y(_05753_),
    .A(net1756),
    .B(\add_result[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11856_ (.B1(_05753_),
    .VDD(VPWR),
    .Y(_01021_),
    .VSS(VGND),
    .A1(net1756),
    .A2(_05752_));
 sg13g2_nand2b_1 _11857_ (.Y(_05754_),
    .B(_05537_),
    .A_N(_05665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11858_ (.Y(_05755_),
    .A(_05536_),
    .B(_05665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11859_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05754_),
    .A2(_05755_),
    .Y(_05756_),
    .B1(\fp16_sum_pipe.seg_reg1.q[21] ));
 sg13g2_inv_1 _11860_ (.VDD(VPWR),
    .Y(_05757_),
    .A(_05497_),
    .VSS(VGND));
 sg13g2_a21oi_1 _11861_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05757_),
    .A2(_05636_),
    .Y(_05758_),
    .B1(net1758));
 sg13g2_o21ai_1 _11862_ (.B1(_05758_),
    .VDD(VPWR),
    .Y(_05759_),
    .VSS(VGND),
    .A1(_05636_),
    .A2(_05489_));
 sg13g2_nand2b_1 _11863_ (.Y(_05760_),
    .B(_05759_),
    .A_N(_05756_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11864_ (.Y(_05761_),
    .A(_05573_),
    .B(\add_result[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11865_ (.B1(_05761_),
    .VDD(VPWR),
    .Y(_01020_),
    .VSS(VGND),
    .A1(_05760_),
    .A2(_05572_));
 sg13g2_nand2_1 _11866_ (.Y(_05762_),
    .A(net1756),
    .B(\add_result[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11867_ (.B1(_05762_),
    .VDD(VPWR),
    .Y(_01019_),
    .VSS(VGND),
    .A1(net1756),
    .A2(_05551_));
 sg13g2_mux2_1 _11868_ (.A0(\add_result[5] ),
    .A1(_05515_),
    .S(net1850),
    .X(_01018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11869_ (.A0(\add_result[4] ),
    .A1(_05481_),
    .S(net1850),
    .X(_01017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11870_ (.A(net1850),
    .B(\add_result[3] ),
    .Y(_05763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11871_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05562_),
    .A2(net1850),
    .Y(_01016_),
    .B1(_05763_));
 sg13g2_mux2_1 _11872_ (.A0(\add_result[2] ),
    .A1(_05568_),
    .S(net1850),
    .X(_01015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11873_ (.A0(\add_result[1] ),
    .A1(_05555_),
    .S(net1850),
    .X(_01014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11874_ (.VDD(VPWR),
    .Y(_05764_),
    .A(\add_result[0] ),
    .VSS(VGND));
 sg13g2_nand3_1 _11875_ (.B(\fp16_sum_pipe.reg3en.q[0] ),
    .C(_05524_),
    .A(_05540_),
    .Y(_05765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11876_ (.B1(_05765_),
    .VDD(VPWR),
    .Y(_01013_),
    .VSS(VGND),
    .A1(net1850),
    .A2(_05764_));
 sg13g2_nor2_1 _11877_ (.A(\fpdiv.reg1en.q[0] ),
    .B(\fpdiv.divider0.state ),
    .Y(_05766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11878_ (.Y(_05767_),
    .A(_05766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11879_ (.Y(_05768_),
    .A(\fpdiv.divider0.counter[1] ),
    .B(\fpdiv.divider0.counter[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11880_ (.A(_02645_),
    .B(_05768_),
    .Y(_05769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11881_ (.Y(_05770_),
    .A(_02644_),
    .B(_05769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11882_ (.Y(_05771_),
    .A(net1718),
    .B(_05770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11883_ (.B1(_05771_),
    .VDD(VPWR),
    .Y(_01012_),
    .VSS(VGND),
    .A1(_02644_),
    .A2(_05767_));
 sg13g2_o21ai_1 _11884_ (.B1(_05767_),
    .VDD(VPWR),
    .Y(_05772_),
    .VSS(VGND),
    .A1(_05769_),
    .A2(_02654_));
 sg13g2_o21ai_1 _11885_ (.B1(_02645_),
    .VDD(VPWR),
    .Y(_05773_),
    .VSS(VGND),
    .A1(_05768_),
    .A2(_02654_));
 sg13g2_and2_1 _11886_ (.A(_05772_),
    .B(_05773_),
    .X(_01011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11887_ (.VDD(VPWR),
    .Y(_05774_),
    .A(\fpdiv.divider0.counter[1] ),
    .VSS(VGND));
 sg13g2_nand3_1 _11888_ (.B(\fpdiv.divider0.state ),
    .C(_05768_),
    .A(_02647_),
    .Y(_05775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11889_ (.B1(_05775_),
    .VDD(VPWR),
    .Y(_01010_),
    .VSS(VGND),
    .A1(_05774_),
    .A2(_05767_));
 sg13g2_nor2_1 _11890_ (.A(\fpdiv.divider0.counter[0] ),
    .B(net1718),
    .Y(_05776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11891_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fpdiv.divider0.counter[0] ),
    .A2(_05767_),
    .Y(_01009_),
    .B1(_05776_));
 sg13g2_xnor2_1 _11892_ (.Y(_05777_),
    .A(\fpmul.reg_a_out[15] ),
    .B(\fpmul.reg_b_out[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11893_ (.A(\fpmul.result[15] ),
    .B(net1876),
    .Y(_05778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05777_),
    .A2(net1876),
    .Y(_01008_),
    .B1(_05778_));
 sg13g2_mux2_1 _11895_ (.A0(\fpmul.seg_reg0.q[53] ),
    .A1(\fpmul.reg_a_out[14] ),
    .S(net1878),
    .X(_01007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11896_ (.A0(\fpmul.seg_reg0.q[52] ),
    .A1(\fpmul.reg_a_out[13] ),
    .S(net1878),
    .X(_01006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11897_ (.A0(\fpmul.seg_reg0.q[51] ),
    .A1(\fpmul.reg_a_out[12] ),
    .S(net1878),
    .X(_01005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11898_ (.VDD(VPWR),
    .Y(_05779_),
    .A(\fpmul.seg_reg0.q[50] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11899_ (.Y(_05780_),
    .A(net1877),
    .B(\fpmul.reg_a_out[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11900_ (.B1(_05780_),
    .VDD(VPWR),
    .Y(_01004_),
    .VSS(VGND),
    .A1(net1877),
    .A2(_05779_));
 sg13g2_mux2_1 _11901_ (.A0(\fpmul.seg_reg0.q[49] ),
    .A1(\fpmul.reg_a_out[10] ),
    .S(net1876),
    .X(_01003_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11902_ (.A0(\fpmul.seg_reg0.q[48] ),
    .A1(\fpmul.reg_a_out[9] ),
    .S(net1876),
    .X(_01002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11903_ (.A0(\fpmul.seg_reg0.q[47] ),
    .A1(\fpmul.reg_a_out[8] ),
    .S(net1876),
    .X(_01001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11904_ (.A0(\fpmul.seg_reg0.q[46] ),
    .A1(\fpmul.reg_a_out[7] ),
    .S(net1876),
    .X(_01000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _11905_ (.A0(\fpmul.seg_reg0.q[45] ),
    .A1(net1854),
    .S(net1880),
    .X(_00999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _11906_ (.Y(_05781_),
    .A(\fpmul.reg_a_out[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11907_ (.A(net1880),
    .B(\fpmul.seg_reg0.q[44] ),
    .Y(_05782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1880),
    .A2(_05781_),
    .Y(_00998_),
    .B1(_05782_));
 sg13g2_inv_2 _11909_ (.Y(_05783_),
    .A(\fpmul.reg_a_out[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11910_ (.A(net1880),
    .B(\fpmul.seg_reg0.q[43] ),
    .Y(_05784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11911_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1880),
    .A2(_05783_),
    .Y(_00997_),
    .B1(_05784_));
 sg13g2_inv_2 _11912_ (.Y(_05785_),
    .A(\fpmul.reg_a_out[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11913_ (.A(net1881),
    .B(\fpmul.seg_reg0.q[42] ),
    .Y(_05786_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11914_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1881),
    .A2(_05785_),
    .Y(_00996_),
    .B1(_05786_));
 sg13g2_inv_1 _11915_ (.VDD(VPWR),
    .Y(_05787_),
    .A(\fpmul.seg_reg0.q[41] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11916_ (.Y(_05788_),
    .A(net1882),
    .B(\fpmul.reg_a_out[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11917_ (.B1(_05788_),
    .VDD(VPWR),
    .Y(_00995_),
    .VSS(VGND),
    .A1(net1881),
    .A2(_05787_));
 sg13g2_inv_1 _11918_ (.VDD(VPWR),
    .Y(_05789_),
    .A(\fpmul.seg_reg0.q[40] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11919_ (.Y(_05790_),
    .A(net1882),
    .B(\fpmul.reg_a_out[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11920_ (.B1(_05790_),
    .VDD(VPWR),
    .Y(_00994_),
    .VSS(VGND),
    .A1(net1881),
    .A2(_05789_));
 sg13g2_inv_1 _11921_ (.VDD(VPWR),
    .Y(_05791_),
    .A(\fpmul.seg_reg0.q[39] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11922_ (.Y(_05792_),
    .A(net1882),
    .B(\fpmul.reg_a_out[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11923_ (.B1(_05792_),
    .VDD(VPWR),
    .Y(_00993_),
    .VSS(VGND),
    .A1(net1882),
    .A2(_05791_));
 sg13g2_inv_1 _11924_ (.VDD(VPWR),
    .Y(_05793_),
    .A(\fpmul.seg_reg0.q[38] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11925_ (.Y(_05794_),
    .A(net1879),
    .B(\fpmul.reg_b_out[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11926_ (.B1(_05794_),
    .VDD(VPWR),
    .Y(_00992_),
    .VSS(VGND),
    .A1(net1879),
    .A2(_05793_));
 sg13g2_inv_1 _11927_ (.VDD(VPWR),
    .Y(_05795_),
    .A(\fpmul.seg_reg0.q[37] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11928_ (.Y(_05796_),
    .A(net1879),
    .B(\fpmul.reg_b_out[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11929_ (.B1(_05796_),
    .VDD(VPWR),
    .Y(_00991_),
    .VSS(VGND),
    .A1(net1879),
    .A2(_05795_));
 sg13g2_inv_1 _11930_ (.VDD(VPWR),
    .Y(_05797_),
    .A(\fpmul.seg_reg0.q[36] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11931_ (.Y(_05798_),
    .A(net1879),
    .B(\fpmul.reg_b_out[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11932_ (.B1(_05798_),
    .VDD(VPWR),
    .Y(_00990_),
    .VSS(VGND),
    .A1(net1879),
    .A2(_05797_));
 sg13g2_inv_1 _11933_ (.VDD(VPWR),
    .Y(_05799_),
    .A(\fpmul.seg_reg0.q[35] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11934_ (.Y(_05800_),
    .A(net1879),
    .B(\fpmul.reg_b_out[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11935_ (.B1(_05800_),
    .VDD(VPWR),
    .Y(_00989_),
    .VSS(VGND),
    .A1(net1879),
    .A2(_05799_));
 sg13g2_inv_1 _11936_ (.VDD(VPWR),
    .Y(_05801_),
    .A(\fpmul.seg_reg0.q[34] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11937_ (.Y(_05802_),
    .A(net1877),
    .B(\fpmul.reg_b_out[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11938_ (.B1(_05802_),
    .VDD(VPWR),
    .Y(_00988_),
    .VSS(VGND),
    .A1(net1874),
    .A2(_05801_));
 sg13g2_inv_1 _11939_ (.VDD(VPWR),
    .Y(_05803_),
    .A(\fpmul.seg_reg0.q[33] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11940_ (.Y(_05804_),
    .A(net1877),
    .B(\fpmul.reg_b_out[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11941_ (.B1(_05804_),
    .VDD(VPWR),
    .Y(_00987_),
    .VSS(VGND),
    .A1(net1874),
    .A2(_05803_));
 sg13g2_inv_1 _11942_ (.VDD(VPWR),
    .Y(_05805_),
    .A(\fpmul.seg_reg0.q[32] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11943_ (.Y(_05806_),
    .A(net1874),
    .B(\fpmul.reg_b_out[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11944_ (.B1(_05806_),
    .VDD(VPWR),
    .Y(_00986_),
    .VSS(VGND),
    .A1(net1874),
    .A2(_05805_));
 sg13g2_inv_1 _11945_ (.VDD(VPWR),
    .Y(_05807_),
    .A(\fpmul.seg_reg0.q[31] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11946_ (.Y(_05808_),
    .A(net1874),
    .B(\fpmul.reg_b_out[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11947_ (.B1(_05808_),
    .VDD(VPWR),
    .Y(_00985_),
    .VSS(VGND),
    .A1(net1874),
    .A2(_05807_));
 sg13g2_inv_1 _11948_ (.VDD(VPWR),
    .Y(_05809_),
    .A(\fpmul.seg_reg0.q[30] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11949_ (.Y(_05810_),
    .A(net1884),
    .B(net1863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11950_ (.B1(_05810_),
    .VDD(VPWR),
    .Y(_00984_),
    .VSS(VGND),
    .A1(net1884),
    .A2(_05809_));
 sg13g2_inv_1 _11951_ (.VDD(VPWR),
    .Y(_05811_),
    .A(\fpmul.seg_reg0.q[29] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11952_ (.Y(_05812_),
    .A(net1883),
    .B(\fpmul.reg_b_out[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11953_ (.B1(_05812_),
    .VDD(VPWR),
    .Y(_00983_),
    .VSS(VGND),
    .A1(net1883),
    .A2(_05811_));
 sg13g2_inv_1 _11954_ (.VDD(VPWR),
    .Y(_05813_),
    .A(\fpmul.seg_reg0.q[28] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11955_ (.Y(_05814_),
    .A(net1882),
    .B(\fpmul.reg_b_out[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11956_ (.B1(_05814_),
    .VDD(VPWR),
    .Y(_00982_),
    .VSS(VGND),
    .A1(net1883),
    .A2(_05813_));
 sg13g2_inv_1 _11957_ (.VDD(VPWR),
    .Y(_05815_),
    .A(\fpmul.seg_reg0.q[27] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11958_ (.Y(_05816_),
    .A(net1883),
    .B(\fpmul.reg_b_out[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11959_ (.B1(_05816_),
    .VDD(VPWR),
    .Y(_00981_),
    .VSS(VGND),
    .A1(net1884),
    .A2(_05815_));
 sg13g2_inv_1 _11960_ (.VDD(VPWR),
    .Y(_05817_),
    .A(\fpmul.seg_reg0.q[26] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11961_ (.Y(_05818_),
    .A(net1884),
    .B(\fpmul.reg_b_out[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11962_ (.B1(_05818_),
    .VDD(VPWR),
    .Y(_00980_),
    .VSS(VGND),
    .A1(net1884),
    .A2(_05817_));
 sg13g2_inv_1 _11963_ (.VDD(VPWR),
    .Y(_05819_),
    .A(\fpmul.seg_reg0.q[25] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11964_ (.Y(_05820_),
    .A(net1883),
    .B(\fpmul.reg_b_out[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11965_ (.B1(_05820_),
    .VDD(VPWR),
    .Y(_00979_),
    .VSS(VGND),
    .A1(net1883),
    .A2(_05819_));
 sg13g2_inv_1 _11966_ (.VDD(VPWR),
    .Y(_05821_),
    .A(\fpmul.seg_reg0.q[24] ),
    .VSS(VGND));
 sg13g2_nand2_1 _11967_ (.Y(_05822_),
    .A(net1884),
    .B(\fpmul.reg_b_out[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11968_ (.B1(_05822_),
    .VDD(VPWR),
    .Y(_00978_),
    .VSS(VGND),
    .A1(net1884),
    .A2(_05821_));
 sg13g2_nand2_1 _11969_ (.Y(_05823_),
    .A(\fpmul.reg_a_out[13] ),
    .B(\fpmul.reg_b_out[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11970_ (.Y(_05824_),
    .A(\fpmul.reg_a_out[14] ),
    .B(\fpmul.reg_b_out[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _11971_ (.B(_05824_),
    .A(_05823_),
    .X(_05825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _11972_ (.B(\fpmul.reg_b_out[12] ),
    .A(\fpmul.reg_a_out[12] ),
    .X(_05826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11973_ (.VDD(VPWR),
    .Y(_05827_),
    .A(_05826_),
    .VSS(VGND));
 sg13g2_nand2_1 _11974_ (.Y(_05828_),
    .A(\fpmul.reg_a_out[11] ),
    .B(\fpmul.reg_b_out[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _11975_ (.B(\fpmul.reg_b_out[11] ),
    .A(\fpmul.reg_a_out[11] ),
    .X(_05829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11976_ (.VDD(VPWR),
    .Y(_05830_),
    .A(_05829_),
    .VSS(VGND));
 sg13g2_nand2_1 _11977_ (.Y(_05831_),
    .A(\fpmul.reg_a_out[10] ),
    .B(\fpmul.reg_b_out[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11978_ (.Y(_05832_),
    .A(\fpmul.reg_a_out[9] ),
    .B(\fpmul.reg_b_out[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11979_ (.VDD(VPWR),
    .Y(_05833_),
    .A(_05832_),
    .VSS(VGND));
 sg13g2_xor2_1 _11980_ (.B(\fpmul.reg_b_out[10] ),
    .A(\fpmul.reg_a_out[10] ),
    .X(_05834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11981_ (.Y(_05835_),
    .A(_05832_),
    .B(_05834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11982_ (.VDD(VPWR),
    .Y(_05836_),
    .A(_05835_),
    .VSS(VGND));
 sg13g2_nand2_1 _11983_ (.Y(_05837_),
    .A(\fpmul.reg_a_out[8] ),
    .B(\fpmul.reg_b_out[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _11984_ (.B(\fpmul.reg_b_out[9] ),
    .A(\fpmul.reg_a_out[9] ),
    .X(_05838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11985_ (.Y(_05839_),
    .A(_05837_),
    .B(_05838_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _11986_ (.A(\fpmul.reg_a_out[7] ),
    .B(\fpmul.reg_b_out[7] ),
    .Y(_05840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _11987_ (.B(\fpmul.reg_b_out[8] ),
    .A(\fpmul.reg_a_out[8] ),
    .X(_05841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _11988_ (.VDD(VPWR),
    .Y(_05842_),
    .A(_05841_),
    .VSS(VGND));
 sg13g2_nor2_1 _11989_ (.A(_05840_),
    .B(_05842_),
    .Y(_05843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _11990_ (.A(_05837_),
    .B_N(_05838_),
    .Y(_05844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _11991_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05839_),
    .A2(_05843_),
    .Y(_05845_),
    .B1(_05844_));
 sg13g2_nor2_1 _11992_ (.A(_05836_),
    .B(_05845_),
    .Y(_05846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _11993_ (.A2(_05834_),
    .A1(_05833_),
    .B1(_05846_),
    .X(_05847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _11994_ (.Y(_05848_),
    .A(_05831_),
    .B(_05829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11995_ (.Y(_05849_),
    .A(_05847_),
    .B(_05848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11996_ (.B1(_05849_),
    .VDD(VPWR),
    .Y(_05850_),
    .VSS(VGND),
    .A1(_05830_),
    .A2(_05831_));
 sg13g2_xnor2_1 _11997_ (.Y(_05851_),
    .A(_05828_),
    .B(_05826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _11998_ (.Y(_05852_),
    .A(_05850_),
    .B(_05851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _11999_ (.B1(_05852_),
    .VDD(VPWR),
    .Y(_05853_),
    .VSS(VGND),
    .A1(_05827_),
    .A2(_05828_));
 sg13g2_nand2_1 _12000_ (.Y(_05854_),
    .A(\fpmul.reg_a_out[12] ),
    .B(\fpmul.reg_b_out[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12001_ (.B(\fpmul.reg_b_out[13] ),
    .A(\fpmul.reg_a_out[13] ),
    .X(_05855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12002_ (.Y(_05856_),
    .A(_05854_),
    .B(_05855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12003_ (.A(_05854_),
    .B_N(_05855_),
    .Y(_05857_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12004_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05853_),
    .A2(_05856_),
    .Y(_05858_),
    .B1(_05857_));
 sg13g2_xnor2_1 _12005_ (.Y(_05859_),
    .A(_05825_),
    .B(_05858_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12006_ (.A(net1875),
    .B(\fpmul.seg_reg0.q[23] ),
    .Y(_05860_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12007_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05859_),
    .A2(net1875),
    .Y(_00977_),
    .B1(_05860_));
 sg13g2_xnor2_1 _12008_ (.Y(_05861_),
    .A(_05856_),
    .B(_05853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12009_ (.A(net1875),
    .B(\fpmul.seg_reg0.q[22] ),
    .Y(_05862_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12010_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05861_),
    .A2(net1875),
    .Y(_00976_),
    .B1(_05862_));
 sg13g2_inv_2 _12011_ (.Y(_05863_),
    .A(\fpmul.seg_reg0.q[21] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12012_ (.A(_05851_),
    .B(_05850_),
    .Y(_05864_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _12013_ (.B(net1878),
    .C(_05852_),
    .Y(_05865_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05864_));
 sg13g2_o21ai_1 _12014_ (.B1(_05865_),
    .VDD(VPWR),
    .Y(_00975_),
    .VSS(VGND),
    .A1(net1877),
    .A2(_05863_));
 sg13g2_xnor2_1 _12015_ (.Y(_05866_),
    .A(_05848_),
    .B(_05847_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12016_ (.A(net1874),
    .B(\fpmul.seg_reg0.q[20] ),
    .Y(_05867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12017_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05866_),
    .A2(net1877),
    .Y(_00974_),
    .B1(_05867_));
 sg13g2_inv_1 _12018_ (.VDD(VPWR),
    .Y(_05868_),
    .A(\fpmul.seg_reg0.q[19] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12019_ (.Y(_05869_),
    .A(_05845_),
    .B(_05836_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _12020_ (.B(net1875),
    .C(_05869_),
    .Y(_05870_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05846_));
 sg13g2_o21ai_1 _12021_ (.B1(_05870_),
    .VDD(VPWR),
    .Y(_00973_),
    .VSS(VGND),
    .A1(net1873),
    .A2(_05868_));
 sg13g2_xnor2_1 _12022_ (.Y(_05871_),
    .A(_05843_),
    .B(_05839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12023_ (.A(net1873),
    .B(\fpmul.seg_reg0.q[18] ),
    .Y(_05872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12024_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05871_),
    .A2(net1873),
    .Y(_00972_),
    .B1(_05872_));
 sg13g2_inv_2 _12025_ (.Y(_05873_),
    .A(\fpmul.seg_reg0.q[17] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12026_ (.Y(_05874_),
    .A(_05842_),
    .B(_05840_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _12027_ (.B(net1873),
    .C(_05874_),
    .Y(_05875_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_05843_));
 sg13g2_o21ai_1 _12028_ (.B1(_05875_),
    .VDD(VPWR),
    .Y(_00971_),
    .VSS(VGND),
    .A1(net1873),
    .A2(_05873_));
 sg13g2_inv_2 _12029_ (.Y(_05876_),
    .A(\fpmul.reg1en.q[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12030_ (.VDD(VPWR),
    .Y(_05877_),
    .A(\fpmul.seg_reg0.q[16] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12031_ (.Y(_05878_),
    .A(\fpmul.reg_a_out[7] ),
    .B(\fpmul.reg_b_out[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12032_ (.A(_05876_),
    .B(_05840_),
    .Y(_05879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12033_ (.Y(_00970_),
    .B1(_05878_),
    .B2(_05879_),
    .A2(_05877_),
    .A1(_05876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12034_ (.Y(_05880_),
    .A(\fpmul.reg_a_out[2] ),
    .B(net1863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12035_ (.VDD(VPWR),
    .Y(_05881_),
    .A(\fpmul.reg_a_out[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12036_ (.Y(_05882_),
    .A(_05880_),
    .B(_05881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12037_ (.B(net1859),
    .C(net1863),
    .A(net1858),
    .Y(_05883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12038_ (.Y(_05884_),
    .A(_05882_),
    .B(_05883_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12039_ (.Y(_05885_),
    .A(net1857),
    .B(net1864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12040_ (.Y(_05886_),
    .A(_05884_),
    .B(_05885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12041_ (.VDD(VPWR),
    .Y(_05887_),
    .A(_05885_),
    .VSS(VGND));
 sg13g2_nand3_1 _12042_ (.B(_05883_),
    .C(_05887_),
    .A(_05882_),
    .Y(_05888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12043_ (.Y(_05889_),
    .A(_05886_),
    .B(_05888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12044_ (.Y(_05890_),
    .A(net1859),
    .B(net1863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _12045_ (.Y(_05891_),
    .A(net1860),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12046_ (.Y(_05892_),
    .A(_05890_),
    .B(_05891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12047_ (.Y(_05893_),
    .A(net1858),
    .B(\fpmul.reg_b_out[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12048_ (.VDD(VPWR),
    .Y(_05894_),
    .A(_05893_),
    .VSS(VGND));
 sg13g2_nand3_1 _12049_ (.B(net1860),
    .C(net1863),
    .A(net1859),
    .Y(_05895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12050_ (.VDD(VPWR),
    .Y(_05896_),
    .A(_05895_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12051_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05892_),
    .A2(_05894_),
    .Y(_05897_),
    .B1(_05896_));
 sg13g2_nand2_1 _12052_ (.Y(_05898_),
    .A(_05889_),
    .B(_05897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12053_ (.Y(_05899_),
    .A(net1855),
    .B(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12054_ (.Y(_05900_),
    .A(net1856),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12055_ (.Y(_05901_),
    .A(net1855),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12056_ (.Y(_05902_),
    .A(net1856),
    .B(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12057_ (.Y(_05903_),
    .A(_05901_),
    .B(_05902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12058_ (.B1(_05903_),
    .VDD(VPWR),
    .Y(_05904_),
    .VSS(VGND),
    .A1(_05899_),
    .A2(_05900_));
 sg13g2_xnor2_1 _12059_ (.Y(_05905_),
    .A(\fpmul.reg_b_out[1] ),
    .B(_05904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12060_ (.A(_05897_),
    .B(_05889_),
    .Y(_05906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12061_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05898_),
    .A2(_05905_),
    .Y(_05907_),
    .B1(_05906_));
 sg13g2_inv_1 _12062_ (.VDD(VPWR),
    .Y(_05908_),
    .A(_05907_),
    .VSS(VGND));
 sg13g2_inv_1 _12063_ (.VDD(VPWR),
    .Y(_05909_),
    .A(_05883_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12064_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05882_),
    .A2(_05887_),
    .Y(_05910_),
    .B1(_05909_));
 sg13g2_inv_1 _12065_ (.VDD(VPWR),
    .Y(_05911_),
    .A(_05910_),
    .VSS(VGND));
 sg13g2_nand2_1 _12066_ (.Y(_05912_),
    .A(\fpmul.reg_a_out[3] ),
    .B(\fpmul.reg_b_out[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12067_ (.VDD(VPWR),
    .Y(_05913_),
    .A(\fpmul.reg_a_out[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12068_ (.Y(_05914_),
    .A(_05912_),
    .B(_05913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12069_ (.B(\fpmul.reg_a_out[2] ),
    .C(net1863),
    .A(net1857),
    .Y(_05915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12070_ (.Y(_05916_),
    .A(net1856),
    .B(net1864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12071_ (.VDD(VPWR),
    .Y(_05917_),
    .A(_05916_),
    .VSS(VGND));
 sg13g2_nand3_1 _12072_ (.B(_05915_),
    .C(_05917_),
    .A(_05914_),
    .Y(_05918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12073_ (.Y(_05919_),
    .A(_05914_),
    .B(_05915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12074_ (.Y(_05920_),
    .A(_05919_),
    .B(_05916_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12075_ (.B(_05918_),
    .C(_05920_),
    .A(_05911_),
    .Y(_05921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12076_ (.Y(_05922_),
    .A(_05920_),
    .B(_05918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12077_ (.Y(_05923_),
    .A(_05922_),
    .B(_05910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12078_ (.Y(_05924_),
    .A(_05921_),
    .B(_05923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12079_ (.Y(_05925_),
    .A(\fpmul.reg_a_out[6] ),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12080_ (.B(_05899_),
    .A(_05925_),
    .X(_05926_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12081_ (.VDD(VPWR),
    .Y(_05927_),
    .A(_05926_),
    .VSS(VGND));
 sg13g2_nand2_1 _12082_ (.Y(_05928_),
    .A(_05924_),
    .B(_05927_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12083_ (.B(_05923_),
    .C(_05926_),
    .A(_05921_),
    .Y(_05929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12084_ (.B(_05928_),
    .C(_05929_),
    .A(_05908_),
    .Y(_05930_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12085_ (.Y(_05931_),
    .A(_05928_),
    .B(_05929_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12086_ (.Y(_05932_),
    .A(_05931_),
    .B(_05907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12087_ (.Y(_05933_),
    .A(_05930_),
    .B(_05932_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12088_ (.A(_05899_),
    .B(_05900_),
    .Y(_05934_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12089_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05903_),
    .A2(net1868),
    .Y(_05935_),
    .B1(_05934_));
 sg13g2_xnor2_1 _12090_ (.Y(_05936_),
    .A(net1867),
    .B(_05935_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12091_ (.VDD(VPWR),
    .Y(_05937_),
    .A(_05936_),
    .VSS(VGND));
 sg13g2_nand2_1 _12092_ (.Y(_05938_),
    .A(_05933_),
    .B(_05937_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12093_ (.B(_05932_),
    .C(_05936_),
    .A(_05930_),
    .Y(_05939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12094_ (.Y(_05940_),
    .A(_05938_),
    .B(_05939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12095_ (.VDD(VPWR),
    .Y(_05941_),
    .A(_05897_),
    .VSS(VGND));
 sg13g2_nand3_1 _12096_ (.B(_05888_),
    .C(_05886_),
    .A(_05941_),
    .Y(_05942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12097_ (.Y(_05943_),
    .A(_05942_),
    .B(_05898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12098_ (.VDD(VPWR),
    .Y(_05944_),
    .A(_05905_),
    .VSS(VGND));
 sg13g2_nand2_1 _12099_ (.Y(_05945_),
    .A(_05943_),
    .B(_05944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12100_ (.B(_05898_),
    .C(_05905_),
    .A(_05942_),
    .Y(_05946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12101_ (.Y(_05947_),
    .A(_05945_),
    .B(_05946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12102_ (.Y(_05948_),
    .A(_05892_),
    .B(_05895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12103_ (.Y(_05949_),
    .A(_05948_),
    .B(_05893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12104_ (.B(_05895_),
    .C(_05894_),
    .A(_05892_),
    .Y(_05950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12105_ (.Y(_05951_),
    .A(_05949_),
    .B(_05950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12106_ (.VDD(VPWR),
    .Y(_05952_),
    .A(_05890_),
    .VSS(VGND));
 sg13g2_nand2_1 _12107_ (.Y(_05953_),
    .A(net1860),
    .B(\fpmul.reg_b_out[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12108_ (.VDD(VPWR),
    .Y(_05954_),
    .A(_05953_),
    .VSS(VGND));
 sg13g2_nand2_1 _12109_ (.Y(_05955_),
    .A(_05952_),
    .B(_05954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12110_ (.Y(_05956_),
    .A(_05951_),
    .B(_05955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12111_ (.Y(_05957_),
    .A(\fpmul.reg_a_out[6] ),
    .B(net1868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12112_ (.VDD(VPWR),
    .Y(_05958_),
    .A(_05957_),
    .VSS(VGND));
 sg13g2_nand2_1 _12113_ (.Y(_05959_),
    .A(net1857),
    .B(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12114_ (.Y(_05960_),
    .A(_05900_),
    .B(_05959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12115_ (.Y(_05961_),
    .A(_05958_),
    .B(_05960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _12116_ (.B(net1858),
    .C(net1860),
    .A(_05952_),
    .Y(_05962_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\fpmul.reg_b_out[5] ));
 sg13g2_inv_1 _12117_ (.VDD(VPWR),
    .Y(_05963_),
    .A(_05962_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12118_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05956_),
    .A2(_05961_),
    .Y(_05964_),
    .B1(_05963_));
 sg13g2_nand2_1 _12119_ (.Y(_05965_),
    .A(_05947_),
    .B(_05964_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12120_ (.Y(_05966_),
    .A(\fpmul.reg_a_out[6] ),
    .B(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12121_ (.Y(_05967_),
    .A(net1857),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12122_ (.A(_05902_),
    .B(_05967_),
    .Y(_05968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12123_ (.A(_05957_),
    .B(_05960_),
    .Y(_05969_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12124_ (.A(_05968_),
    .B(_05969_),
    .Y(_05970_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12125_ (.B(_05970_),
    .A(_05966_),
    .X(_05971_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12126_ (.A(_05964_),
    .B(_05947_),
    .Y(_05972_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05965_),
    .A2(_05971_),
    .Y(_05973_),
    .B1(_05972_));
 sg13g2_nand2_1 _12128_ (.Y(_05974_),
    .A(_05940_),
    .B(_05973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12129_ (.A(_05966_),
    .B(_05970_),
    .Y(_05975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12130_ (.A(_05973_),
    .B(_05940_),
    .Y(_05976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12131_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05974_),
    .A2(_05975_),
    .Y(_05977_),
    .B1(_05976_));
 sg13g2_inv_1 _12132_ (.VDD(VPWR),
    .Y(_05978_),
    .A(_05977_),
    .VSS(VGND));
 sg13g2_nor2_1 _12133_ (.A(_05907_),
    .B(_05931_),
    .Y(_05979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12134_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05932_),
    .A2(_05936_),
    .Y(_05980_),
    .B1(_05979_));
 sg13g2_inv_1 _12135_ (.VDD(VPWR),
    .Y(_05981_),
    .A(_05980_),
    .VSS(VGND));
 sg13g2_nand2_1 _12136_ (.Y(_05982_),
    .A(\fpmul.reg_a_out[6] ),
    .B(\fpmul.reg_b_out[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12137_ (.A(_05982_),
    .B(_05901_),
    .Y(_05983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12138_ (.A(_05910_),
    .B(_05922_),
    .Y(_05984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12139_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05923_),
    .A2(_05926_),
    .Y(_05985_),
    .B1(_05984_));
 sg13g2_inv_1 _12140_ (.VDD(VPWR),
    .Y(_05986_),
    .A(_05985_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12141_ (.Y(_05987_),
    .A(net1866),
    .B(_05982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12142_ (.VDD(VPWR),
    .Y(_05988_),
    .A(_05915_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12143_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05914_),
    .A2(_05917_),
    .Y(_05989_),
    .B1(_05988_));
 sg13g2_inv_1 _12144_ (.VDD(VPWR),
    .Y(_05990_),
    .A(_05989_),
    .VSS(VGND));
 sg13g2_nand2_1 _12145_ (.Y(_05991_),
    .A(net1856),
    .B(\fpmul.reg_b_out[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12146_ (.Y(_05992_),
    .A(_05991_),
    .B(_05785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12147_ (.B(\fpmul.reg_a_out[3] ),
    .C(\fpmul.reg_b_out[6] ),
    .A(net1856),
    .Y(_05993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12148_ (.Y(_05994_),
    .A(_05992_),
    .B(_05993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12149_ (.Y(_05995_),
    .A(net1855),
    .B(net1864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12150_ (.Y(_05996_),
    .A(_05994_),
    .B(_05995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12151_ (.VDD(VPWR),
    .Y(_05997_),
    .A(_05995_),
    .VSS(VGND));
 sg13g2_nand3_1 _12152_ (.B(_05993_),
    .C(_05997_),
    .A(_05992_),
    .Y(_05998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12153_ (.B(_05996_),
    .C(_05998_),
    .A(_05990_),
    .Y(_05999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12154_ (.Y(_06000_),
    .A(_05996_),
    .B(_05998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12155_ (.Y(_06001_),
    .A(_06000_),
    .B(_05989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12156_ (.Y(_06002_),
    .A(_05999_),
    .B(_06001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12157_ (.Y(_06003_),
    .B(_06002_),
    .A_N(_05987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12158_ (.B(_06001_),
    .C(_05987_),
    .A(_05999_),
    .Y(_06004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12159_ (.B(_06003_),
    .C(_06004_),
    .A(_05986_),
    .Y(_06005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12160_ (.Y(_06006_),
    .A(_06003_),
    .B(_06004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12161_ (.Y(_06007_),
    .A(_06006_),
    .B(_05985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12162_ (.Y(_06008_),
    .A(_06005_),
    .B(_06007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12163_ (.Y(_06009_),
    .B(_06008_),
    .A_N(_05983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12164_ (.B(_06007_),
    .C(_05983_),
    .A(_06005_),
    .Y(_06010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12165_ (.B(_06009_),
    .C(_06010_),
    .A(_05981_),
    .Y(_06011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12166_ (.Y(_06012_),
    .A(_06009_),
    .B(_06010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12167_ (.Y(_06013_),
    .A(_06012_),
    .B(_05980_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12168_ (.Y(_06014_),
    .A(_06011_),
    .B(_06013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _12169_ (.Y(_06015_),
    .A(\fpmul.reg_b_out[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12170_ (.A(_06015_),
    .B(_05935_),
    .Y(_06016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12171_ (.VDD(VPWR),
    .Y(_06017_),
    .A(_06016_),
    .VSS(VGND));
 sg13g2_nand2_1 _12172_ (.Y(_06018_),
    .A(_06014_),
    .B(_06017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12173_ (.B(_06013_),
    .C(_06016_),
    .A(_06011_),
    .Y(_06019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12174_ (.B(_06018_),
    .C(_06019_),
    .A(_05978_),
    .Y(_06020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_72_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_72_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12176_ (.VDD(VPWR),
    .Y(_06022_),
    .A(_06005_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12177_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06007_),
    .A2(_05983_),
    .Y(_06023_),
    .B1(_06022_));
 sg13g2_inv_1 _12178_ (.VDD(VPWR),
    .Y(_06024_),
    .A(_06023_),
    .VSS(VGND));
 sg13g2_inv_2 _12179_ (.Y(_06025_),
    .A(\fpmul.reg_b_out[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12180_ (.A(_06025_),
    .B(_05925_),
    .Y(_06026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _12181_ (.A(_05998_),
    .B(_05993_),
    .X(_06027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12182_ (.VDD(VPWR),
    .Y(_06028_),
    .A(_06027_),
    .VSS(VGND));
 sg13g2_nand2_1 _12183_ (.Y(_06029_),
    .A(\fpmul.reg_a_out[6] ),
    .B(net1864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12184_ (.VDD(VPWR),
    .Y(_06030_),
    .A(_06029_),
    .VSS(VGND));
 sg13g2_inv_1 _12185_ (.VDD(VPWR),
    .Y(_06031_),
    .A(\fpmul.reg_b_out[6] ),
    .VSS(VGND));
 sg13g2_o21ai_1 _12186_ (.B1(_05783_),
    .VDD(VPWR),
    .Y(_06032_),
    .VSS(VGND),
    .A1(_05781_),
    .A2(_06031_));
 sg13g2_inv_1 _12187_ (.VDD(VPWR),
    .Y(_06033_),
    .A(_05991_),
    .VSS(VGND));
 sg13g2_nand2_1 _12188_ (.Y(_06034_),
    .A(_06033_),
    .B(net1855),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12189_ (.Y(_06035_),
    .A(_06032_),
    .B(_06034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12190_ (.Y(_06036_),
    .A(_06030_),
    .B(_06035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12191_ (.Y(_06037_),
    .A(_06028_),
    .B(_06036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12192_ (.Y(_06038_),
    .A(_06029_),
    .B(_06035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12193_ (.Y(_06039_),
    .A(_06038_),
    .B(_06027_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12194_ (.Y(_06040_),
    .A(_06037_),
    .B(_06039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12195_ (.Y(_06041_),
    .A(_06040_),
    .B(_06025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12196_ (.B(_06039_),
    .C(\fpmul.reg_b_out[4] ),
    .A(_06037_),
    .Y(_06042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12197_ (.Y(_06043_),
    .A(_06041_),
    .B(_06042_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12198_ (.VDD(VPWR),
    .Y(_06044_),
    .A(_05999_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12199_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06001_),
    .A2(_05987_),
    .Y(_06045_),
    .B1(_06044_));
 sg13g2_nand2_1 _12200_ (.Y(_06046_),
    .A(_06043_),
    .B(_06045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12201_ (.VDD(VPWR),
    .Y(_06047_),
    .A(_06045_),
    .VSS(VGND));
 sg13g2_nand3_1 _12202_ (.B(_06042_),
    .C(_06047_),
    .A(_06041_),
    .Y(_06048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12203_ (.Y(_06049_),
    .A(_06046_),
    .B(_06048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12204_ (.Y(_06050_),
    .B(_06049_),
    .A_N(_06026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12205_ (.B(_06048_),
    .C(_06026_),
    .A(_06046_),
    .Y(_06051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12206_ (.Y(_06052_),
    .A(_06050_),
    .B(_06051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12207_ (.Y(_06053_),
    .A(_06024_),
    .B(_06052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12208_ (.VDD(VPWR),
    .Y(_06054_),
    .A(_06011_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12209_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06013_),
    .A2(_06016_),
    .Y(_06055_),
    .B1(_06054_));
 sg13g2_xnor2_1 _12210_ (.Y(_06056_),
    .A(_06053_),
    .B(_06055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12211_ (.VDD(VPWR),
    .Y(_06057_),
    .A(_06056_),
    .VSS(VGND));
 sg13g2_nand2b_1 _12212_ (.Y(_06058_),
    .B(_06053_),
    .A_N(_06055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12213_ (.B1(_06058_),
    .VDD(VPWR),
    .Y(_06059_),
    .VSS(VGND),
    .A1(_06020_),
    .A2(_06057_));
 sg13g2_nand2_1 _12214_ (.Y(_06060_),
    .A(_06018_),
    .B(_06019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12215_ (.Y(_06061_),
    .A(_06060_),
    .B(_05977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12216_ (.B(_06020_),
    .C(_06061_),
    .A(_06056_),
    .Y(_06062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12217_ (.Y(_06063_),
    .A(net1856),
    .B(net1868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12218_ (.Y(_06064_),
    .A(net1858),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12219_ (.Y(_06065_),
    .A(net1859),
    .B(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12220_ (.Y(_06066_),
    .A(_06064_),
    .B(_06065_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12221_ (.Y(_06067_),
    .A(_06063_),
    .B(_06066_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12222_ (.A(_05953_),
    .B(_06067_),
    .Y(_06068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12223_ (.Y(_06069_),
    .A(net1860),
    .B(net1863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12224_ (.Y(_06070_),
    .A(net1859),
    .B(\fpmul.reg_b_out[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12225_ (.B(_06070_),
    .A(_06069_),
    .X(_06071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12226_ (.Y(_06072_),
    .A(net1855),
    .B(net1868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12227_ (.Y(_06073_),
    .A(net1858),
    .B(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12228_ (.Y(_06074_),
    .A(_05967_),
    .B(_06073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12229_ (.Y(_06075_),
    .A(_06072_),
    .B(_06074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12230_ (.B(_06075_),
    .A(_06071_),
    .X(_06076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12231_ (.Y(_06077_),
    .A(_06068_),
    .B(_06076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12232_ (.Y(_06078_),
    .A(\fpmul.reg_a_out[6] ),
    .B(net1869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12233_ (.Y(_06079_),
    .A(net1856),
    .B(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12234_ (.Y(_06080_),
    .A(net1859),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12235_ (.A(_06073_),
    .B(_06080_),
    .Y(_06081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12236_ (.A(_06063_),
    .B(_06066_),
    .Y(_06082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12237_ (.A(_06081_),
    .B(_06082_),
    .Y(_06083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12238_ (.B(_06083_),
    .A(_06079_),
    .X(_06084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12239_ (.Y(_06085_),
    .A(_06078_),
    .B(_06084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12240_ (.Y(_06086_),
    .A(_06077_),
    .B(_06085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12241_ (.Y(_06087_),
    .B(_06068_),
    .A_N(_06076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12242_ (.Y(_06088_),
    .A(_06086_),
    .B(_06087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12243_ (.Y(_06089_),
    .A(net1855),
    .B(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12244_ (.A(_05959_),
    .B(_06064_),
    .Y(_06090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12245_ (.A(_06072_),
    .B(_06074_),
    .Y(_06091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _12246_ (.A(_06090_),
    .B(_06091_),
    .Y(_06092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12247_ (.Y(_06093_),
    .A(_06089_),
    .B(_06092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12248_ (.Y(_06094_),
    .A(net1869),
    .B(_06093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12249_ (.Y(_06095_),
    .A(_05956_),
    .B(_05962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12250_ (.Y(_06096_),
    .B(_06095_),
    .A_N(_05961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12251_ (.B(_05962_),
    .C(_05961_),
    .A(_05956_),
    .Y(_06097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12252_ (.Y(_06098_),
    .A(_06096_),
    .B(_06097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12253_ (.A(_06075_),
    .B_N(_06071_),
    .Y(_06099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12254_ (.VDD(VPWR),
    .Y(_06100_),
    .A(_06099_),
    .VSS(VGND));
 sg13g2_nand2_1 _12255_ (.Y(_06101_),
    .A(_06098_),
    .B(_06100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12256_ (.B(_06097_),
    .C(_06099_),
    .A(_06096_),
    .Y(_06102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12257_ (.Y(_06103_),
    .A(_06101_),
    .B(_06102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12258_ (.Y(_06104_),
    .B(_06103_),
    .A_N(_06094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12259_ (.B(_06094_),
    .C(_06102_),
    .A(_06101_),
    .Y(_06105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12260_ (.Y(_06106_),
    .A(_06104_),
    .B(_06105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12261_ (.Y(_06107_),
    .B(_06106_),
    .A_N(_06088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12262_ (.VDD(VPWR),
    .Y(_06108_),
    .A(_06078_),
    .VSS(VGND));
 sg13g2_nor2_1 _12263_ (.A(_06079_),
    .B(_06083_),
    .Y(_06109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12264_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06084_),
    .A2(_06108_),
    .Y(_06110_),
    .B1(_06109_));
 sg13g2_inv_1 _12265_ (.VDD(VPWR),
    .Y(_06111_),
    .A(_06110_),
    .VSS(VGND));
 sg13g2_nand3_1 _12266_ (.B(_06104_),
    .C(_06105_),
    .A(_06088_),
    .Y(_06112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12267_ (.VDD(VPWR),
    .Y(_06113_),
    .A(_06112_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12268_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06107_),
    .A2(_06111_),
    .Y(_06114_),
    .B1(_06113_));
 sg13g2_inv_1 _12269_ (.VDD(VPWR),
    .Y(_06115_),
    .A(_06102_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12270_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06101_),
    .A2(_06094_),
    .Y(_06116_),
    .B1(_06115_));
 sg13g2_inv_1 _12271_ (.VDD(VPWR),
    .Y(_06117_),
    .A(_06116_),
    .VSS(VGND));
 sg13g2_inv_1 _12272_ (.VDD(VPWR),
    .Y(_06118_),
    .A(_05964_),
    .VSS(VGND));
 sg13g2_nand3_1 _12273_ (.B(_05946_),
    .C(_05945_),
    .A(_06118_),
    .Y(_06119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12274_ (.Y(_06120_),
    .A(_06119_),
    .B(_05965_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12275_ (.VDD(VPWR),
    .Y(_06121_),
    .A(_05971_),
    .VSS(VGND));
 sg13g2_nand2_1 _12276_ (.Y(_06122_),
    .A(_06120_),
    .B(_06121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12277_ (.B(_05965_),
    .C(_05971_),
    .A(_06119_),
    .Y(_06123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12278_ (.B(_06122_),
    .C(_06123_),
    .A(_06117_),
    .Y(_06124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12279_ (.Y(_06125_),
    .A(_06122_),
    .B(_06123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12280_ (.Y(_06126_),
    .A(_06125_),
    .B(_06116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12281_ (.Y(_06127_),
    .A(_06124_),
    .B(_06126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12282_ (.Y(_06128_),
    .A(_06092_),
    .B(_06089_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12283_ (.A(_06089_),
    .B(_06092_),
    .Y(_06129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12284_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06128_),
    .A2(net1869),
    .Y(_06130_),
    .B1(_06129_));
 sg13g2_nand2_1 _12285_ (.Y(_06131_),
    .A(_06127_),
    .B(_06130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12286_ (.VDD(VPWR),
    .Y(_06132_),
    .A(_06130_),
    .VSS(VGND));
 sg13g2_nand3_1 _12287_ (.B(_06126_),
    .C(_06132_),
    .A(_06124_),
    .Y(_06133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12288_ (.Y(_06134_),
    .A(_06131_),
    .B(_06133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12289_ (.A(_06114_),
    .B(_06134_),
    .Y(_06135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12290_ (.VDD(VPWR),
    .Y(_06136_),
    .A(_05973_),
    .VSS(VGND));
 sg13g2_nand3_1 _12291_ (.B(_05939_),
    .C(_05938_),
    .A(_06136_),
    .Y(_06137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12292_ (.Y(_06138_),
    .A(_06137_),
    .B(_05974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12293_ (.Y(_06139_),
    .B(_06138_),
    .A_N(_05975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12294_ (.B(_05974_),
    .C(_05975_),
    .A(_06137_),
    .Y(_06140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12295_ (.Y(_06141_),
    .A(_06139_),
    .B(_06140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12296_ (.VDD(VPWR),
    .Y(_06142_),
    .A(_06124_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12297_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06126_),
    .A2(_06132_),
    .Y(_06143_),
    .B1(_06142_));
 sg13g2_nand2_1 _12298_ (.Y(_06144_),
    .A(_06141_),
    .B(_06143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12299_ (.A(_06143_),
    .B(_06141_),
    .Y(_06145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12300_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06135_),
    .A2(_06144_),
    .Y(_06146_),
    .B1(_06145_));
 sg13g2_nor2_1 _12301_ (.A(_06062_),
    .B(_06146_),
    .Y(_06147_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12302_ (.A(_06059_),
    .B(_06147_),
    .Y(_06148_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12303_ (.B(_06141_),
    .A(_06143_),
    .X(_06149_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12304_ (.VDD(VPWR),
    .Y(_06150_),
    .A(_06114_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12305_ (.Y(_06151_),
    .A(_06150_),
    .B(_06134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12306_ (.Y(_06152_),
    .A(_06149_),
    .B(_06151_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12307_ (.A(_06062_),
    .B(_06152_),
    .Y(_06153_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12308_ (.VDD(VPWR),
    .Y(_06154_),
    .A(_06077_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12309_ (.Y(_06155_),
    .A(_06108_),
    .B(_06084_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12310_ (.Y(_06156_),
    .A(_06154_),
    .B(_06155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12311_ (.Y(_06157_),
    .A(_06156_),
    .B(_06086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12312_ (.Y(_06158_),
    .A(_05954_),
    .B(_06067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12313_ (.Y(_06159_),
    .A(net1855),
    .B(net1869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12314_ (.Y(_06160_),
    .A(net1857),
    .B(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12315_ (.Y(_06161_),
    .A(net1860),
    .B(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12316_ (.Y(_06162_),
    .A(_06080_),
    .B(_06161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12317_ (.Y(_06163_),
    .A(net1857),
    .B(net1868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12318_ (.VDD(VPWR),
    .Y(_06164_),
    .A(_06163_),
    .VSS(VGND));
 sg13g2_nand2_2 _12319_ (.Y(_06165_),
    .A(net1860),
    .B(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12320_ (.A(_06065_),
    .B(_06165_),
    .Y(_06166_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _12321_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_06166_),
    .Y(_06167_),
    .A2(_06164_),
    .A1(_06162_));
 sg13g2_xor2_1 _12322_ (.B(_06167_),
    .A(_06160_),
    .X(_06168_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12323_ (.Y(_06169_),
    .B(_06168_),
    .A_N(_06159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12324_ (.Y(_06170_),
    .A(_06160_),
    .B(_06167_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12325_ (.Y(_06171_),
    .A(_06170_),
    .B(_06159_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12326_ (.B(_06169_),
    .C(_06171_),
    .A(_06158_),
    .Y(_06172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout119 (.A(net128),
    .X(net119),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12328_ (.Y(_06174_),
    .A(_06157_),
    .B(_06172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12329_ (.A(_06160_),
    .B(_06167_),
    .Y(_06175_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12330_ (.A(_06175_),
    .B_N(_06169_),
    .Y(_06176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12331_ (.VDD(VPWR),
    .Y(_06177_),
    .A(_06176_),
    .VSS(VGND));
 sg13g2_inv_1 _12332_ (.VDD(VPWR),
    .Y(_06178_),
    .A(_06172_),
    .VSS(VGND));
 sg13g2_nand3_1 _12333_ (.B(_06086_),
    .C(_06178_),
    .A(_06156_),
    .Y(_06179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12334_ (.VDD(VPWR),
    .Y(_06180_),
    .A(_06179_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12335_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06174_),
    .A2(_06177_),
    .Y(_06181_),
    .B1(_06180_));
 sg13g2_nand2_1 _12336_ (.Y(_06182_),
    .A(_06107_),
    .B(_06112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12337_ (.Y(_06183_),
    .A(_06182_),
    .B(_06110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12338_ (.B(_06112_),
    .C(_06111_),
    .A(_06107_),
    .Y(_06184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _12339_ (.B(_06183_),
    .C(_06184_),
    .Y(_06185_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06181_));
 sg13g2_nand2_1 _12340_ (.Y(_06186_),
    .A(_06174_),
    .B(_06179_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12341_ (.Y(_06187_),
    .A(_06186_),
    .B(_06176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12342_ (.B(_06179_),
    .C(_06177_),
    .A(_06174_),
    .Y(_06188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12343_ (.Y(_06189_),
    .A(net1856),
    .B(net1869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12344_ (.VDD(VPWR),
    .Y(_06190_),
    .A(_06189_),
    .VSS(VGND));
 sg13g2_nand2_1 _12345_ (.Y(_06191_),
    .A(net1858),
    .B(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12346_ (.Y(_06192_),
    .A(net1858),
    .B(net1868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12347_ (.A(_06165_),
    .B(_06192_),
    .Y(_06193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12348_ (.Y(_06194_),
    .A(_06191_),
    .B(_06193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12349_ (.Y(_06195_),
    .A(_06190_),
    .B(_06194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12350_ (.B1(_06162_),
    .VDD(VPWR),
    .Y(_06196_),
    .VSS(VGND),
    .A1(_06065_),
    .A2(_06165_));
 sg13g2_xnor2_1 _12351_ (.Y(_06197_),
    .A(_06164_),
    .B(_06196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12352_ (.A(_06195_),
    .B_N(_06197_),
    .Y(_06198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12353_ (.Y(_06199_),
    .A(_06169_),
    .B(_06171_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12354_ (.Y(_06200_),
    .B(_06199_),
    .A_N(_06158_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12355_ (.Y(_06201_),
    .A(_06200_),
    .B(_06172_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12356_ (.Y(_06202_),
    .B(_06201_),
    .A_N(_06198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _12357_ (.A(_06015_),
    .B(_06165_),
    .C(_06192_),
    .Y(_06203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _12358_ (.A2(_06190_),
    .A1(_06194_),
    .B1(_06203_),
    .X(_06204_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12359_ (.B(_06172_),
    .C(_06198_),
    .A(_06200_),
    .Y(_06205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12360_ (.VDD(VPWR),
    .Y(_06206_),
    .A(_06205_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12361_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06202_),
    .A2(_06204_),
    .Y(_06207_),
    .B1(_06206_));
 sg13g2_inv_1 _12362_ (.VDD(VPWR),
    .Y(_06208_),
    .A(_06207_),
    .VSS(VGND));
 sg13g2_nand3_1 _12363_ (.B(_06188_),
    .C(_06208_),
    .A(_06187_),
    .Y(_06209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12364_ (.Y(_06210_),
    .A(_06185_),
    .B(_06209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12365_ (.Y(_06211_),
    .A(_06202_),
    .B(_06205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12366_ (.B(_06211_),
    .A(_06204_),
    .X(_06212_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12367_ (.B(_06192_),
    .A(_06165_),
    .X(_06213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12368_ (.Y(_06214_),
    .A(net1857),
    .B(net1869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12369_ (.Y(_06215_),
    .A(net1859),
    .B(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12370_ (.B(_06215_),
    .A(_06214_),
    .X(_06216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12371_ (.Y(_06217_),
    .A(_06213_),
    .B(_06216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12372_ (.B(_06195_),
    .A(_06197_),
    .X(_06218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12373_ (.A(_06217_),
    .B(_06218_),
    .Y(_06219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _12374_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_06220_),
    .B(_06215_),
    .A(_06214_));
 sg13g2_xnor2_1 _12375_ (.Y(_06221_),
    .A(_06217_),
    .B(_06218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12376_ (.A(_06220_),
    .B(_06221_),
    .Y(_06222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12377_ (.A(_06219_),
    .B(_06222_),
    .Y(_06223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12378_ (.Y(_06224_),
    .A(_06212_),
    .B(_06223_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12379_ (.Y(_06225_),
    .A(net1858),
    .B(\fpmul.reg_b_out[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12380_ (.B1(_06225_),
    .VDD(VPWR),
    .Y(_06226_),
    .VSS(VGND),
    .A1(_05891_),
    .A2(_06015_));
 sg13g2_nand2_1 _12381_ (.Y(_06227_),
    .A(net1859),
    .B(\fpmul.reg_b_out[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12382_ (.VDD(VPWR),
    .Y(_06228_),
    .A(_06227_),
    .VSS(VGND));
 sg13g2_nor3_1 _12383_ (.A(_05891_),
    .B(_06015_),
    .C(_06225_),
    .Y(_06229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12384_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06226_),
    .A2(_06228_),
    .Y(_06230_),
    .B1(_06229_));
 sg13g2_xor2_1 _12385_ (.B(_06216_),
    .A(_06213_),
    .X(_06231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12386_ (.VDD(VPWR),
    .Y(_06232_),
    .A(_06231_),
    .VSS(VGND));
 sg13g2_nor2_2 _12387_ (.A(_06230_),
    .B(_06232_),
    .Y(_06233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12388_ (.VDD(VPWR),
    .Y(_06234_),
    .A(_06233_),
    .VSS(VGND));
 sg13g2_inv_1 _12389_ (.VDD(VPWR),
    .Y(_06235_),
    .A(_06229_),
    .VSS(VGND));
 sg13g2_nand3_1 _12390_ (.B(net1860),
    .C(\fpmul.reg_b_out[0] ),
    .A(_06228_),
    .Y(_06236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _12391_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_06230_),
    .C1(_06236_),
    .B1(_06232_),
    .A1(_06235_),
    .Y(_06237_),
    .A2(_06226_));
 sg13g2_inv_1 _12392_ (.VDD(VPWR),
    .Y(_06238_),
    .A(_06237_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12393_ (.Y(_06239_),
    .A(_06220_),
    .B(_06221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06234_),
    .A2(_06238_),
    .Y(_06240_),
    .B1(_06239_));
 sg13g2_nor2_1 _12395_ (.A(_06223_),
    .B(_06212_),
    .Y(_06241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12396_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06224_),
    .A2(_06240_),
    .Y(_06242_),
    .B1(_06241_));
 sg13g2_nand2_1 _12397_ (.Y(_06243_),
    .A(_06187_),
    .B(_06188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12398_ (.Y(_06244_),
    .A(_06243_),
    .B(_06207_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12399_ (.Y(_06245_),
    .A(_06244_),
    .B(_06209_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12400_ (.A(_06242_),
    .B(_06245_),
    .Y(_06246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12401_ (.A(_06210_),
    .B(_06246_),
    .Y(_06247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12402_ (.Y(_06248_),
    .A(_06183_),
    .B(_06184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12403_ (.Y(_06249_),
    .A(_06248_),
    .B(_06181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _12404_ (.A(_06247_),
    .B_N(_06249_),
    .Y(_06250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12405_ (.Y(_06251_),
    .A(_06153_),
    .B(_06250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12406_ (.Y(_06252_),
    .A(_06148_),
    .B(_06251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12407_ (.B(_06051_),
    .C(_06024_),
    .A(_06050_),
    .Y(_06253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12408_ (.Y(_06254_),
    .A(net1854),
    .B(\fpmul.reg_b_out[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12409_ (.Y(_06255_),
    .A(_05781_),
    .B(_06254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12410_ (.Y(_06256_),
    .A(net1864),
    .B(_06255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12411_ (.Y(_06257_),
    .B1(_06030_),
    .B2(_06032_),
    .A2(_06033_),
    .A1(net1855),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12412_ (.B(_06257_),
    .A(_06256_),
    .X(_06258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _12413_ (.A(_06042_),
    .B(_06037_),
    .X(_06259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12414_ (.Y(_06260_),
    .A(_06258_),
    .B(_06259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _12415_ (.A(_06051_),
    .B(_06048_),
    .X(_06261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12417_ (.Y(_06263_),
    .A(_06260_),
    .B(_06261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12418_ (.B(_06263_),
    .A(_06253_),
    .X(_06264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12419_ (.VDD(VPWR),
    .Y(_06265_),
    .A(_06264_),
    .VSS(VGND));
 sg13g2_nor2_1 _12420_ (.A(net1854),
    .B(\fpmul.reg_b_out[6] ),
    .Y(_06266_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12421_ (.VDD(VPWR),
    .Y(_06267_),
    .A(_06254_),
    .VSS(VGND));
 sg13g2_nor2_1 _12422_ (.A(_06266_),
    .B(_06267_),
    .Y(_06268_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12423_ (.Y(_06269_),
    .B(net1864),
    .A_N(_06255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12424_ (.VDD(VPWR),
    .Y(_06270_),
    .A(_06266_),
    .VSS(VGND));
 sg13g2_o21ai_1 _12425_ (.B1(_06270_),
    .VDD(VPWR),
    .Y(_06271_),
    .VSS(VGND),
    .A1(\fpmul.reg_a_out[5] ),
    .A2(_06254_));
 sg13g2_nor2b_1 _12426_ (.A(_06257_),
    .B_N(_06256_),
    .Y(_06272_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _12427_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_06271_),
    .C1(_06272_),
    .B1(_06269_),
    .A1(_05997_),
    .Y(_06273_),
    .A2(_06268_));
 sg13g2_nor2_1 _12428_ (.A(_06258_),
    .B(_06259_),
    .Y(_06274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12429_ (.Y(_06275_),
    .A(_06273_),
    .B(_06274_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12430_ (.A(_06260_),
    .B(_06261_),
    .Y(_06276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12431_ (.Y(_06277_),
    .A(_06275_),
    .B(_06276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12432_ (.A(_06265_),
    .B_N(_06277_),
    .Y(_06278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12433_ (.Y(_06279_),
    .A(_06252_),
    .B(_06278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12434_ (.A(_06253_),
    .B(_06263_),
    .Y(_06280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _12435_ (.A(_06275_),
    .B(_06260_),
    .C(_06261_),
    .Y(_06281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06277_),
    .A2(_06280_),
    .Y(_06282_),
    .B1(_06281_));
 sg13g2_nand2_1 _12437_ (.Y(_06283_),
    .A(_06279_),
    .B(_06282_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12438_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06270_),
    .A2(_05997_),
    .Y(_06284_),
    .B1(_06267_));
 sg13g2_nor2b_1 _12439_ (.A(_06272_),
    .B_N(_06284_),
    .Y(_06285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12440_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06267_),
    .A2(_06272_),
    .Y(_06286_),
    .B1(_06285_));
 sg13g2_and2_1 _12441_ (.A(_06274_),
    .B(_06273_),
    .X(_06287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12442_ (.Y(_06288_),
    .A(_06286_),
    .B(_06287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12443_ (.Y(_06289_),
    .A(_06283_),
    .B(_06288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12444_ (.Y(_06290_),
    .B(_06287_),
    .A_N(_06286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12445_ (.B(_06285_),
    .C(_06290_),
    .A(_06289_),
    .Y(_06291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12446_ (.Y(_06292_),
    .A(_06291_),
    .B(net1870),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12447_ (.Y(_06293_),
    .A(_05876_),
    .B(\fpmul.seg_reg0.q[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12448_ (.Y(_00969_),
    .A(_06292_),
    .B(_06293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12449_ (.A(_06288_),
    .B(_06283_),
    .Y(_06294_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _12450_ (.B(net1870),
    .C(_06289_),
    .Y(_06295_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06294_));
 sg13g2_nand2_1 _12451_ (.Y(_06296_),
    .A(_05876_),
    .B(\fpmul.seg_reg0.q[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12452_ (.Y(_00968_),
    .A(_06295_),
    .B(_06296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12453_ (.Y(_06297_),
    .A(_06252_),
    .B(_06264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12454_ (.Y(_06298_),
    .B(_06297_),
    .A_N(_06280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12455_ (.Y(_06299_),
    .A(_06277_),
    .B(_06298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12456_ (.A(net1870),
    .B(\fpmul.seg_reg0.q[13] ),
    .Y(_06300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12457_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06299_),
    .A2(net1870),
    .Y(_00967_),
    .B1(_06300_));
 sg13g2_inv_1 _12458_ (.VDD(VPWR),
    .Y(_06301_),
    .A(\fpmul.seg_reg0.q[12] ),
    .VSS(VGND));
 sg13g2_nand3_1 _12459_ (.B(_06251_),
    .C(_06265_),
    .A(_06148_),
    .Y(_06302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12460_ (.B(_06302_),
    .C(net1870),
    .A(_06297_),
    .Y(_06303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12461_ (.B1(_06303_),
    .VDD(VPWR),
    .Y(_00966_),
    .VSS(VGND),
    .A1(net1870),
    .A2(_06301_));
 sg13g2_inv_1 _12462_ (.VDD(VPWR),
    .Y(_06304_),
    .A(\fpmul.seg_reg0.q[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12463_ (.Y(_06305_),
    .A(_06020_),
    .B(_06061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12464_ (.Y(_06306_),
    .B(_06250_),
    .A_N(_06152_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12465_ (.Y(_06307_),
    .A(_06306_),
    .B(_06146_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12466_ (.Y(_06308_),
    .B(_06307_),
    .A_N(_06305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12467_ (.Y(_06309_),
    .A(_06308_),
    .B(_06020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12468_ (.Y(_06310_),
    .A(_06309_),
    .B(_06056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12469_ (.B(_06020_),
    .C(_06057_),
    .A(_06308_),
    .Y(_06311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12470_ (.B(_06311_),
    .C(net1870),
    .A(_06310_),
    .Y(_06312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12471_ (.B1(_06312_),
    .VDD(VPWR),
    .Y(_00965_),
    .VSS(VGND),
    .A1(net1871),
    .A2(_06304_));
 sg13g2_inv_1 _12472_ (.VDD(VPWR),
    .Y(_06313_),
    .A(\fpmul.seg_reg0.q[10] ),
    .VSS(VGND));
 sg13g2_nand3_1 _12473_ (.B(_06305_),
    .C(_06146_),
    .A(_06306_),
    .Y(_06314_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12474_ (.B(_06314_),
    .C(net1871),
    .A(_06308_),
    .Y(_06315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12475_ (.B1(_06315_),
    .VDD(VPWR),
    .Y(_00964_),
    .VSS(VGND),
    .A1(net1871),
    .A2(_06313_));
 sg13g2_a21oi_1 _12476_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06250_),
    .A2(_06151_),
    .Y(_06316_),
    .B1(_06135_));
 sg13g2_xor2_1 _12477_ (.B(_06316_),
    .A(_06149_),
    .X(_06317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12478_ (.A(net1872),
    .B(\fpmul.seg_reg0.q[9] ),
    .Y(_06318_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12479_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06317_),
    .A2(net1872),
    .Y(_00963_),
    .B1(_06318_));
 sg13g2_xnor2_1 _12480_ (.Y(_06319_),
    .A(_06151_),
    .B(_06250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12481_ (.A(net1872),
    .B(\fpmul.seg_reg0.q[8] ),
    .Y(_06320_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12482_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06319_),
    .A2(net1872),
    .Y(_00962_),
    .B1(_06320_));
 sg13g2_nand2_1 _12483_ (.Y(_06321_),
    .A(_06185_),
    .B(_06249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12484_ (.A(_06246_),
    .B_N(_06209_),
    .Y(_06322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12485_ (.Y(_06323_),
    .A(_06321_),
    .B(_06322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12486_ (.A(net1872),
    .B(\fpmul.seg_reg0.q[7] ),
    .Y(_06324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12487_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06323_),
    .A2(net1872),
    .Y(_00961_),
    .B1(_06324_));
 sg13g2_xnor2_1 _12488_ (.Y(_06325_),
    .A(_06242_),
    .B(_06245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12489_ (.A(net1872),
    .B(\fpmul.seg_reg0.q[6] ),
    .Y(_06326_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12490_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06325_),
    .A2(net1872),
    .Y(_00960_),
    .B1(_06326_));
 sg13g2_nor2b_1 _12491_ (.A(_06241_),
    .B_N(_06224_),
    .Y(_06327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12492_ (.Y(_06328_),
    .A(_06240_),
    .B(_06327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12493_ (.A(net1871),
    .B(\fpmul.seg_reg0.q[5] ),
    .Y(_06329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12494_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06328_),
    .A2(net1871),
    .Y(_00959_),
    .B1(_06329_));
 sg13g2_nor2_1 _12495_ (.A(_06233_),
    .B(_06238_),
    .Y(_06330_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12496_ (.Y(_06331_),
    .A(_06233_),
    .B(_06239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12497_ (.Y(_06332_),
    .A(_06330_),
    .B(_06331_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12498_ (.A(net1871),
    .B(\fpmul.seg_reg0.q[4] ),
    .Y(_06333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12499_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06332_),
    .A2(net1871),
    .Y(_00958_),
    .B1(_06333_));
 sg13g2_nor2_1 _12500_ (.A(\fpmul.reg_a_out[15] ),
    .B(net1951),
    .Y(_06334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12501_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03327_),
    .A2(net1951),
    .Y(_00957_),
    .B1(_06334_));
 sg13g2_nor2_1 _12502_ (.A(\fpmul.reg_a_out[14] ),
    .B(net1953),
    .Y(_06335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12503_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05357_),
    .A2(net1953),
    .Y(_00956_),
    .B1(_06335_));
 sg13g2_nor2_1 _12504_ (.A(\fpmul.reg_a_out[13] ),
    .B(net1951),
    .Y(_06336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12505_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05359_),
    .A2(net1951),
    .Y(_00955_),
    .B1(_06336_));
 sg13g2_inv_1 _12506_ (.VDD(VPWR),
    .Y(_06337_),
    .A(\acc_sub.x2[12] ),
    .VSS(VGND));
 sg13g2_nor2_1 _12507_ (.A(\fpmul.reg_a_out[12] ),
    .B(net1953),
    .Y(_06338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06337_),
    .A2(net1953),
    .Y(_00954_),
    .B1(_06338_));
 sg13g2_inv_1 _12509_ (.VDD(VPWR),
    .Y(_06339_),
    .A(\acc_sub.x2[11] ),
    .VSS(VGND));
 sg13g2_nor2_1 _12510_ (.A(\fpmul.reg_a_out[11] ),
    .B(net1953),
    .Y(_06340_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12511_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06339_),
    .A2(net1953),
    .Y(_00953_),
    .B1(_06340_));
 sg13g2_inv_1 _12512_ (.VDD(VPWR),
    .Y(_06341_),
    .A(\acc_sub.x2[10] ),
    .VSS(VGND));
 sg13g2_nor2_1 _12513_ (.A(\fpmul.reg_a_out[10] ),
    .B(net1953),
    .Y(_06342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12514_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06341_),
    .A2(net1953),
    .Y(_00952_),
    .B1(_06342_));
 sg13g2_nor2_1 _12515_ (.A(\fpmul.reg_a_out[9] ),
    .B(net1958),
    .Y(_06343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12516_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_05367_),
    .A2(net1958),
    .Y(_00951_),
    .B1(_06343_));
 sg13g2_nor2_1 _12517_ (.A(\fpmul.reg_a_out[8] ),
    .B(net1955),
    .Y(_06344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03601_),
    .A2(net1955),
    .Y(_00950_),
    .B1(_06344_));
 sg13g2_nor2_1 _12519_ (.A(\fpmul.reg_a_out[7] ),
    .B(net1951),
    .Y(_06345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12520_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_03603_),
    .A2(net1951),
    .Y(_00949_),
    .B1(_06345_));
 sg13g2_inv_2 _12521_ (.Y(_06346_),
    .A(\acc_sub.x2[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12522_ (.A(net1854),
    .B(net1959),
    .Y(_06347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12523_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06346_),
    .A2(net1959),
    .Y(_00948_),
    .B1(_06347_));
 sg13g2_nand2_1 _12524_ (.Y(_06348_),
    .A(\acc_sub.x2[5] ),
    .B(net1956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12525_ (.B1(_06348_),
    .VDD(VPWR),
    .Y(_00947_),
    .VSS(VGND),
    .A1(net1956),
    .A2(_05781_));
 sg13g2_nand2_1 _12526_ (.Y(_06349_),
    .A(\acc_sub.x2[4] ),
    .B(net1955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12527_ (.B1(_06349_),
    .VDD(VPWR),
    .Y(_00946_),
    .VSS(VGND),
    .A1(net1956),
    .A2(_05783_));
 sg13g2_nand2_1 _12528_ (.Y(_06350_),
    .A(\acc_sub.x2[3] ),
    .B(net1956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12529_ (.B1(_06350_),
    .VDD(VPWR),
    .Y(_00945_),
    .VSS(VGND),
    .A1(net1956),
    .A2(_05785_));
 sg13g2_nand2_1 _12530_ (.Y(_06351_),
    .A(\acc_sub.x2[2] ),
    .B(net1954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12531_ (.B1(_06351_),
    .VDD(VPWR),
    .Y(_00944_),
    .VSS(VGND),
    .A1(net1954),
    .A2(_05913_));
 sg13g2_nand2_1 _12532_ (.Y(_06352_),
    .A(\acc_sub.x2[1] ),
    .B(net1955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12533_ (.B1(_06352_),
    .VDD(VPWR),
    .Y(_00943_),
    .VSS(VGND),
    .A1(net1954),
    .A2(_05881_));
 sg13g2_nand2_1 _12534_ (.Y(_06353_),
    .A(\acc_sub.x2[0] ),
    .B(net1957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12535_ (.B1(_06353_),
    .VDD(VPWR),
    .Y(_00942_),
    .VSS(VGND),
    .A1(net1957),
    .A2(_05891_));
 sg13g2_buf_2 fanout77 (.A(net80),
    .X(net77),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _12537_ (.A(_02648_),
    .Y(_06354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12538_ (.Y(_06355_),
    .A(_05374_),
    .B(_05376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _12539_ (.B(_05378_),
    .C(_05380_),
    .A(_05372_),
    .Y(_06356_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_02722_));
 sg13g2_nor4_1 _12540_ (.A(\fpdiv.reg_a_out[10] ),
    .B(\fpdiv.reg_a_out[9] ),
    .C(\fpdiv.reg_a_out[8] ),
    .D(\fpdiv.reg_a_out[7] ),
    .Y(_06357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _12541_ (.A(\fpdiv.reg_a_out[14] ),
    .B(\fpdiv.reg_a_out[13] ),
    .C(\fpdiv.reg_a_out[12] ),
    .D(\fpdiv.reg_a_out[11] ),
    .Y(_06358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12542_ (.Y(_06359_),
    .A(_06357_),
    .B(_06358_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_2 _12543_ (.A(\fpdiv.divider0.dividend[5] ),
    .B(_06355_),
    .C(_06356_),
    .Y(_06360_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_06359_));
 sg13g2_nor4_1 _12544_ (.A(\fpdiv.divider0.divisor[6] ),
    .B(\fpdiv.divider0.divisor[5] ),
    .C(\fpdiv.divider0.divisor[4] ),
    .D(\fpdiv.reg_b_out[14] ),
    .Y(_06361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _12545_ (.A(\fpdiv.divider0.divisor[10] ),
    .B(\fpdiv.divider0.divisor[9] ),
    .C(\fpdiv.divider0.divisor[8] ),
    .D(\fpdiv.divider0.divisor[7] ),
    .Y(_06362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12546_ (.Y(_06363_),
    .A(_06361_),
    .B(_06362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _12547_ (.A(\fpdiv.reg_b_out[13] ),
    .B(\fpdiv.reg_b_out[12] ),
    .C(\fpdiv.reg_b_out[11] ),
    .D(\fpdiv.reg_b_out[10] ),
    .Y(_06364_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _12548_ (.B(_05387_),
    .C(_05389_),
    .A(_06364_),
    .Y(_06365_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05391_));
 sg13g2_nor2_1 _12549_ (.A(_06363_),
    .B(_06365_),
    .Y(_06366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout89 (.A(net91),
    .X(net89),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12551_ (.B(\fpdiv.reg_b_out[15] ),
    .A(\fpdiv.reg_a_out[15] ),
    .X(_06368_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12552_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06360_),
    .A2(net1735),
    .Y(_06369_),
    .B1(_06368_));
 sg13g2_nand2_1 _12553_ (.Y(_06370_),
    .A(_06354_),
    .B(\div_result[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12554_ (.B1(_06370_),
    .VDD(VPWR),
    .Y(_00941_),
    .VSS(VGND),
    .A1(_06354_),
    .A2(_06369_));
 sg13g2_inv_1 _12555_ (.VDD(VPWR),
    .Y(_06371_),
    .A(\div_result[14] ),
    .VSS(VGND));
 sg13g2_buf_2 fanout88 (.A(net92),
    .X(net88),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12557_ (.A(\fpdiv.reg_b_out[11] ),
    .B(_05363_),
    .Y(_06373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12558_ (.Y(_06374_),
    .A(\fpdiv.reg_a_out[12] ),
    .B(\fpdiv.reg_b_out[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12559_ (.B(_06374_),
    .A(_06373_),
    .X(_06375_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12560_ (.Y(_06376_),
    .A(\fpdiv.reg_a_out[8] ),
    .B(\fpdiv.reg_b_out[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12561_ (.VDD(VPWR),
    .Y(_06377_),
    .A(_06376_),
    .VSS(VGND));
 sg13g2_nor3_1 _12562_ (.A(_05370_),
    .B(\fpdiv.reg_b_out[7] ),
    .C(_06377_),
    .Y(_06378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12563_ (.Y(_06379_),
    .A(_05389_),
    .B(\fpdiv.reg_a_out[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12564_ (.Y(_06380_),
    .A(\fpdiv.reg_a_out[9] ),
    .B(\fpdiv.reg_b_out[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12565_ (.Y(_06381_),
    .A(_06379_),
    .B(_06380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12566_ (.A(_06379_),
    .B_N(_06380_),
    .Y(_06382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06378_),
    .A2(_06381_),
    .Y(_06383_),
    .B1(_06382_));
 sg13g2_nand2_1 _12568_ (.Y(_06384_),
    .A(_05387_),
    .B(\fpdiv.reg_a_out[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12569_ (.Y(_06385_),
    .A(\fpdiv.reg_a_out[10] ),
    .B(\fpdiv.reg_b_out[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12570_ (.Y(_06386_),
    .A(_06384_),
    .B(_06385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12571_ (.Y(_06387_),
    .B(_06386_),
    .A_N(_06383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12572_ (.Y(_06388_),
    .B(_06385_),
    .A_N(_06384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12573_ (.Y(_06389_),
    .A(_06387_),
    .B(_06388_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12574_ (.A(\fpdiv.reg_b_out[10] ),
    .B(_05365_),
    .Y(_06390_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12575_ (.Y(_06391_),
    .A(\fpdiv.reg_a_out[11] ),
    .B(\fpdiv.reg_b_out[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12576_ (.B(_06391_),
    .A(_06390_),
    .X(_06392_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _12577_ (.A(_06391_),
    .B(_06390_),
    .X(_06393_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _12578_ (.A2(_06392_),
    .A1(_06389_),
    .B1(_06393_),
    .X(_06394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12579_ (.Y(_06395_),
    .A(_06375_),
    .B(_06394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12580_ (.B(_06389_),
    .A(_06392_),
    .X(_06396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12581_ (.B(_06378_),
    .A(_06381_),
    .X(_06397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12582_ (.B1(_06377_),
    .VDD(VPWR),
    .Y(_06398_),
    .VSS(VGND),
    .A1(_05370_),
    .A2(\fpdiv.reg_b_out[7] ));
 sg13g2_nand2b_1 _12583_ (.Y(_06399_),
    .B(_06398_),
    .A_N(_06378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12584_ (.Y(_06400_),
    .A(\fpdiv.reg_a_out[7] ),
    .B(\fpdiv.reg_b_out[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _12585_ (.A(net1852),
    .B(_06400_),
    .Y(_06401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12586_ (.Y(_06402_),
    .A(_06399_),
    .B(_06401_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12587_ (.A(_06397_),
    .B(_06402_),
    .Y(_06403_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12588_ (.VDD(VPWR),
    .Y(_06404_),
    .A(_06403_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12589_ (.Y(_06405_),
    .A(_06386_),
    .B(_06383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12590_ (.A(_06404_),
    .B(_06405_),
    .Y(_06406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _12591_ (.A(_06396_),
    .B_N(_06406_),
    .Y(_06407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12592_ (.Y(_06408_),
    .A(_06395_),
    .B(_06407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12593_ (.A(\fpdiv.reg_b_out[12] ),
    .B(_05361_),
    .Y(_06409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12594_ (.Y(_06410_),
    .A(\fpdiv.reg_a_out[13] ),
    .B(\fpdiv.reg_b_out[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12595_ (.B(_06410_),
    .A(_06409_),
    .X(_06411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _12596_ (.A(_06374_),
    .B(_06373_),
    .X(_06412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _12597_ (.A2(_06375_),
    .A1(_06394_),
    .B1(_06412_),
    .X(_06413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12598_ (.B(_06413_),
    .A(_06411_),
    .X(_06414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12599_ (.B(_06414_),
    .A(_06408_),
    .X(_06415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12600_ (.B(_06395_),
    .A(_06407_),
    .X(_06416_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12601_ (.Y(_06417_),
    .A(_06406_),
    .B(_06396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12602_ (.Y(_06418_),
    .A(_06403_),
    .B(_06405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12603_ (.B(_06402_),
    .A(_06397_),
    .X(_06419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12604_ (.B(_06399_),
    .A(_06401_),
    .X(_06420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _12605_ (.A(net1851),
    .Y(_06421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12606_ (.Y(_06422_),
    .A(_06421_),
    .B(_05348_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12607_ (.B1(_06422_),
    .VDD(VPWR),
    .Y(_06423_),
    .VSS(VGND),
    .A1(_06421_),
    .A2(\fpdiv.div_out[4] ));
 sg13g2_nand2_1 _12608_ (.Y(_06424_),
    .A(\fpdiv.div_out[11] ),
    .B(\fpdiv.div_out[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12609_ (.B1(_06424_),
    .VDD(VPWR),
    .Y(_06425_),
    .VSS(VGND),
    .A1(\fpdiv.div_out[11] ),
    .A2(_05350_));
 sg13g2_buf_2 fanout72 (.A(net2),
    .X(net72),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12611_ (.VDD(VPWR),
    .Y(_06427_),
    .A(_06425_),
    .VSS(VGND));
 sg13g2_nor2_1 _12612_ (.A(_06423_),
    .B(_06427_),
    .Y(_06428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12613_ (.Y(_06429_),
    .A(\fpdiv.div_out[11] ),
    .B(\fpdiv.div_out[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12614_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06421_),
    .A2(\fpdiv.div_out[0] ),
    .Y(_06430_),
    .B1(\fpdiv.div_out[1] ));
 sg13g2_and3_1 _12615_ (.X(_06431_),
    .A(_06425_),
    .B(_06429_),
    .C(_06430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12616_ (.A(_06427_),
    .B(_06431_),
    .Y(_06432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12617_ (.A(_06428_),
    .B(_06432_),
    .Y(_06433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12618_ (.Y(_06434_),
    .A(_05339_),
    .B(net1851),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12619_ (.B1(_06434_),
    .VDD(VPWR),
    .Y(_06435_),
    .VSS(VGND),
    .A1(net1851),
    .A2(\fpdiv.div_out[8] ));
 sg13g2_nand2_1 _12620_ (.Y(_06436_),
    .A(_06421_),
    .B(_05342_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12621_ (.B1(_06436_),
    .VDD(VPWR),
    .Y(_06437_),
    .VSS(VGND),
    .A1(_06421_),
    .A2(\fpdiv.div_out[8] ));
 sg13g2_buf_1 place1743 (.A(net1742),
    .X(net1743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12623_ (.Y(_06439_),
    .A(_05342_),
    .B(net1852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12624_ (.B1(_06439_),
    .VDD(VPWR),
    .Y(_06440_),
    .VSS(VGND),
    .A1(net1852),
    .A2(\fpdiv.div_out[6] ));
 sg13g2_nand2_1 _12625_ (.Y(_06441_),
    .A(_05345_),
    .B(net1852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12626_ (.B1(_06441_),
    .VDD(VPWR),
    .Y(_06442_),
    .VSS(VGND),
    .A1(net1852),
    .A2(\fpdiv.div_out[4] ));
 sg13g2_nor2_1 _12627_ (.A(_06442_),
    .B(_06423_),
    .Y(_06443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12628_ (.Y(_06444_),
    .A(net1852),
    .B(\fpdiv.div_out[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12629_ (.VDD(VPWR),
    .Y(_06445_),
    .A(_06444_),
    .VSS(VGND));
 sg13g2_a21oi_1 _12630_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06421_),
    .A2(\fpdiv.div_out[5] ),
    .Y(_06446_),
    .B1(_06445_));
 sg13g2_inv_1 _12631_ (.VDD(VPWR),
    .Y(_06447_),
    .A(_06446_),
    .VSS(VGND));
 sg13g2_nand2_1 _12632_ (.Y(_06448_),
    .A(_06443_),
    .B(_06447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12633_ (.A(_06440_),
    .B(_06448_),
    .Y(_06449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12634_ (.VDD(VPWR),
    .Y(_06450_),
    .A(_06449_),
    .VSS(VGND));
 sg13g2_nor2_1 _12635_ (.A(_06437_),
    .B(_06450_),
    .Y(_06451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12636_ (.VDD(VPWR),
    .Y(_06452_),
    .A(_06451_),
    .VSS(VGND));
 sg13g2_nor2_1 _12637_ (.A(_06435_),
    .B(_06452_),
    .Y(_06453_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12638_ (.Y(_06454_),
    .A(_06421_),
    .B(_05337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12639_ (.Y(_06455_),
    .A(net1851),
    .B(\fpdiv.div_out[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12640_ (.B1(_06455_),
    .VDD(VPWR),
    .Y(_06456_),
    .VSS(VGND),
    .A1(net1851),
    .A2(_05339_));
 sg13g2_nand3_1 _12641_ (.B(_06454_),
    .C(_06456_),
    .A(_06453_),
    .Y(_06457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12642_ (.VDD(VPWR),
    .Y(_06458_),
    .A(_06457_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12643_ (.Y(_06459_),
    .A(net1852),
    .B(_06400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _12644_ (.B(_06458_),
    .C(_06459_),
    .Y(_06460_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06433_));
 sg13g2_nor2_1 _12645_ (.A(_06420_),
    .B(_06460_),
    .Y(_06461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12646_ (.Y(_06462_),
    .B(_06461_),
    .A_N(_06419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12647_ (.A(_06418_),
    .B(_06462_),
    .Y(_06463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12648_ (.VDD(VPWR),
    .Y(_06464_),
    .A(_06463_),
    .VSS(VGND));
 sg13g2_nor2_1 _12649_ (.A(_06417_),
    .B(_06464_),
    .Y(_06465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12650_ (.VDD(VPWR),
    .Y(_06466_),
    .A(_06465_),
    .VSS(VGND));
 sg13g2_nor2_1 _12651_ (.A(_06416_),
    .B(_06466_),
    .Y(_06467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12652_ (.Y(_06468_),
    .B(_06467_),
    .A_N(_06415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12653_ (.A(_06408_),
    .B(_06414_),
    .Y(_06469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12654_ (.Y(_06470_),
    .A(_05385_),
    .B(\fpdiv.reg_a_out[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12655_ (.Y(_06471_),
    .A(\fpdiv.reg_a_out[14] ),
    .B(\fpdiv.reg_b_out[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12656_ (.B(_06471_),
    .A(_06470_),
    .X(_06472_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _12657_ (.A(_06410_),
    .B(_06409_),
    .X(_06473_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12658_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06413_),
    .A2(_06411_),
    .Y(_06474_),
    .B1(_06473_));
 sg13g2_xnor2_1 _12659_ (.Y(_06475_),
    .A(_06472_),
    .B(_06474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12660_ (.Y(_06476_),
    .A(_06469_),
    .B(_06475_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12661_ (.B(_06476_),
    .A(_06468_),
    .X(_06477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _12662_ (.Y(_06478_),
    .A(_06366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _12663_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_06354_),
    .Y(_06479_),
    .A2(_06360_),
    .A1(_06478_));
 sg13g2_o21ai_1 _12664_ (.B1(_06479_),
    .VDD(VPWR),
    .Y(_06480_),
    .VSS(VGND),
    .A1(net1735),
    .A2(_06477_));
 sg13g2_o21ai_1 _12665_ (.B1(_06480_),
    .VDD(VPWR),
    .Y(_00940_),
    .VSS(VGND),
    .A1(_06371_),
    .A2(net1741));
 sg13g2_inv_2 _12666_ (.Y(_06481_),
    .A(_06479_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12667_ (.Y(_06482_),
    .B(_06415_),
    .A_N(_06467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06468_),
    .A2(_06482_),
    .Y(_06483_),
    .B1(net1735));
 sg13g2_nand2_1 _12669_ (.Y(_06484_),
    .A(_06354_),
    .B(\div_result[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12670_ (.B1(_06484_),
    .VDD(VPWR),
    .Y(_00939_),
    .VSS(VGND),
    .A1(_06481_),
    .A2(_06483_));
 sg13g2_inv_1 _12671_ (.VDD(VPWR),
    .Y(_06485_),
    .A(\div_result[12] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _12672_ (.Y(_06486_),
    .A(_06416_),
    .B(_06465_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12673_ (.B1(_06479_),
    .VDD(VPWR),
    .Y(_06487_),
    .VSS(VGND),
    .A1(net1735),
    .A2(_06486_));
 sg13g2_o21ai_1 _12674_ (.B1(_06487_),
    .VDD(VPWR),
    .Y(_00938_),
    .VSS(VGND),
    .A1(_06485_),
    .A2(net1741));
 sg13g2_inv_1 _12675_ (.VDD(VPWR),
    .Y(_06488_),
    .A(\div_result[11] ),
    .VSS(VGND));
 sg13g2_nor2_1 _12676_ (.A(_06354_),
    .B(net1735),
    .Y(_06489_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12677_ (.VDD(VPWR),
    .Y(_06490_),
    .A(_06360_),
    .VSS(VGND));
 sg13g2_nand2_1 _12678_ (.Y(_06491_),
    .A(_06464_),
    .B(_06417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12679_ (.B(_06490_),
    .C(_06491_),
    .A(_06466_),
    .Y(_06492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12680_ (.Y(_00937_),
    .B1(_06489_),
    .B2(_06492_),
    .A2(_06354_),
    .A1(_06488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12681_ (.Y(_06493_),
    .A(_06462_),
    .B(_06418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12682_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06464_),
    .A2(_06493_),
    .Y(_06494_),
    .B1(net1735));
 sg13g2_nand2_1 _12683_ (.Y(_06495_),
    .A(_06354_),
    .B(\div_result[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12684_ (.B1(_06495_),
    .VDD(VPWR),
    .Y(_00936_),
    .VSS(VGND),
    .A1(_06481_),
    .A2(_06494_));
 sg13g2_inv_1 _12685_ (.VDD(VPWR),
    .Y(_06496_),
    .A(\div_result[9] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _12686_ (.Y(_06497_),
    .A(_06419_),
    .B(_06461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12687_ (.B1(_06479_),
    .VDD(VPWR),
    .Y(_06498_),
    .VSS(VGND),
    .A1(net1735),
    .A2(_06497_));
 sg13g2_o21ai_1 _12688_ (.B1(_06498_),
    .VDD(VPWR),
    .Y(_00935_),
    .VSS(VGND),
    .A1(_06496_),
    .A2(net1741));
 sg13g2_inv_1 _12689_ (.VDD(VPWR),
    .Y(_06499_),
    .A(\div_result[8] ),
    .VSS(VGND));
 sg13g2_xor2_1 _12690_ (.B(_06460_),
    .A(_06420_),
    .X(_06500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12691_ (.B1(_06479_),
    .VDD(VPWR),
    .Y(_06501_),
    .VSS(VGND),
    .A1(net1734),
    .A2(_06500_));
 sg13g2_o21ai_1 _12692_ (.B1(_06501_),
    .VDD(VPWR),
    .Y(_00934_),
    .VSS(VGND),
    .A1(_06499_),
    .A2(net1741));
 sg13g2_inv_1 _12693_ (.VDD(VPWR),
    .Y(_06502_),
    .A(\div_result[7] ),
    .VSS(VGND));
 sg13g2_inv_1 _12694_ (.VDD(VPWR),
    .Y(_06503_),
    .A(_06431_),
    .VSS(VGND));
 sg13g2_inv_1 _12695_ (.VDD(VPWR),
    .Y(_06504_),
    .A(_06432_),
    .VSS(VGND));
 sg13g2_nor2_1 _12696_ (.A(_06435_),
    .B(_06437_),
    .Y(_06505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _12697_ (.B(_06454_),
    .C(_06456_),
    .A(_06449_),
    .Y(_06506_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_06505_));
 sg13g2_a21oi_1 _12698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06503_),
    .A2(_06504_),
    .Y(_06507_),
    .B1(_06506_));
 sg13g2_xor2_1 _12699_ (.B(_06507_),
    .A(_06459_),
    .X(_06508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12700_ (.B1(_06479_),
    .VDD(VPWR),
    .Y(_06509_),
    .VSS(VGND),
    .A1(net1734),
    .A2(_06508_));
 sg13g2_o21ai_1 _12701_ (.B1(_06509_),
    .VDD(VPWR),
    .Y(_00933_),
    .VSS(VGND),
    .A1(_06502_),
    .A2(net1741));
 sg13g2_inv_2 _12702_ (.Y(_06510_),
    .A(\div_result[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12703_ (.Y(_06511_),
    .A(_06453_),
    .B(_06425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12704_ (.Y(_06512_),
    .A(_06456_),
    .B(_06511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _12705_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_06481_),
    .Y(_06513_),
    .A2(_06490_),
    .A1(net1735));
 sg13g2_buf_2 fanout137 (.A(net138),
    .X(net137),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12707_ (.B1(_06513_),
    .VDD(VPWR),
    .Y(_06515_),
    .VSS(VGND),
    .A1(net1734),
    .A2(_06512_));
 sg13g2_o21ai_1 _12708_ (.B1(_06515_),
    .VDD(VPWR),
    .Y(_00932_),
    .VSS(VGND),
    .A1(_06510_),
    .A2(_02648_));
 sg13g2_inv_1 _12709_ (.VDD(VPWR),
    .Y(_06516_),
    .A(\div_result[5] ),
    .VSS(VGND));
 sg13g2_o21ai_1 _12710_ (.B1(_06435_),
    .VDD(VPWR),
    .Y(_06517_),
    .VSS(VGND),
    .A1(_06427_),
    .A2(_06452_));
 sg13g2_a21oi_1 _12711_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06517_),
    .A2(_06511_),
    .Y(_06518_),
    .B1(net1734));
 sg13g2_nand2b_1 _12712_ (.Y(_06519_),
    .B(_06513_),
    .A_N(_06518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12713_ (.B1(_06519_),
    .VDD(VPWR),
    .Y(_00931_),
    .VSS(VGND),
    .A1(_06516_),
    .A2(net1741));
 sg13g2_inv_1 _12714_ (.VDD(VPWR),
    .Y(_06520_),
    .A(\div_result[4] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12715_ (.Y(_06521_),
    .A(_06504_),
    .B(_06423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12716_ (.Y(_06522_),
    .A(_06450_),
    .B(_06437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _12717_ (.B(_06521_),
    .C(_06522_),
    .A(_06452_),
    .Y(_06523_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_06425_));
 sg13g2_nand2b_1 _12718_ (.Y(_06524_),
    .B(_06433_),
    .A_N(_06437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12719_ (.B(_06478_),
    .C(_06524_),
    .A(_06523_),
    .Y(_06525_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12720_ (.Y(_06526_),
    .A(_06525_),
    .B(_06513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12721_ (.B1(_06526_),
    .VDD(VPWR),
    .Y(_00930_),
    .VSS(VGND),
    .A1(_06520_),
    .A2(net1741));
 sg13g2_inv_1 _12722_ (.VDD(VPWR),
    .Y(_06527_),
    .A(\div_result[3] ),
    .VSS(VGND));
 sg13g2_inv_1 _12723_ (.VDD(VPWR),
    .Y(_06528_),
    .A(_06428_),
    .VSS(VGND));
 sg13g2_nor2_1 _12724_ (.A(_06442_),
    .B(_06528_),
    .Y(_06529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12725_ (.Y(_06530_),
    .A(_06529_),
    .B(_06447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _12726_ (.B(_06530_),
    .A(_06440_),
    .X(_06531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12727_ (.B1(_06513_),
    .VDD(VPWR),
    .Y(_06532_),
    .VSS(VGND),
    .A1(net1734),
    .A2(_06531_));
 sg13g2_o21ai_1 _12728_ (.B1(_06532_),
    .VDD(VPWR),
    .Y(_00929_),
    .VSS(VGND),
    .A1(_06527_),
    .A2(_02648_));
 sg13g2_inv_1 _12729_ (.VDD(VPWR),
    .Y(_06533_),
    .A(\div_result[2] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _12730_ (.Y(_06534_),
    .A(_06446_),
    .B(_06529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12731_ (.B1(_06513_),
    .VDD(VPWR),
    .Y(_06535_),
    .VSS(VGND),
    .A1(net1734),
    .A2(_06534_));
 sg13g2_o21ai_1 _12732_ (.B1(_06535_),
    .VDD(VPWR),
    .Y(_00928_),
    .VSS(VGND),
    .A1(_06533_),
    .A2(_02648_));
 sg13g2_inv_1 _12733_ (.VDD(VPWR),
    .Y(_06536_),
    .A(\div_result[1] ),
    .VSS(VGND));
 sg13g2_xnor2_1 _12734_ (.Y(_06537_),
    .A(_06442_),
    .B(_06428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12735_ (.B1(_06513_),
    .VDD(VPWR),
    .Y(_06538_),
    .VSS(VGND),
    .A1(net1734),
    .A2(_06537_));
 sg13g2_o21ai_1 _12736_ (.B1(_06538_),
    .VDD(VPWR),
    .Y(_00927_),
    .VSS(VGND),
    .A1(_06536_),
    .A2(_02648_));
 sg13g2_inv_2 _12737_ (.Y(_06539_),
    .A(\div_result[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12738_ (.B1(_06521_),
    .VDD(VPWR),
    .Y(_06540_),
    .VSS(VGND),
    .A1(_06528_),
    .A2(_06458_));
 sg13g2_o21ai_1 _12739_ (.B1(_06478_),
    .VDD(VPWR),
    .Y(_06541_),
    .VSS(VGND),
    .A1(_06507_),
    .A2(_06540_));
 sg13g2_nand2_1 _12740_ (.Y(_06542_),
    .A(_06541_),
    .B(_06513_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12741_ (.B1(_06542_),
    .VDD(VPWR),
    .Y(_00926_),
    .VSS(VGND),
    .A1(_06539_),
    .A2(_02648_));
 sg13g2_mux2_1 _12742_ (.A0(\fpmul.reg_b_out[15] ),
    .A1(\fp16_res_pipe.x2[15] ),
    .S(net1951),
    .X(_00925_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12743_ (.A0(\fpmul.reg_b_out[14] ),
    .A1(\fp16_res_pipe.x2[14] ),
    .S(net1952),
    .X(_00924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12744_ (.A0(\fpmul.reg_b_out[13] ),
    .A1(\fp16_res_pipe.x2[13] ),
    .S(net1952),
    .X(_00923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12745_ (.A0(\fpmul.reg_b_out[12] ),
    .A1(\fp16_res_pipe.x2[12] ),
    .S(net1952),
    .X(_00922_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12746_ (.A0(\fpmul.reg_b_out[11] ),
    .A1(\fp16_res_pipe.x2[11] ),
    .S(net1952),
    .X(_00921_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12747_ (.A0(\fpmul.reg_b_out[10] ),
    .A1(\fp16_res_pipe.x2[10] ),
    .S(net1952),
    .X(_00920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12748_ (.A0(\fpmul.reg_b_out[9] ),
    .A1(\fp16_res_pipe.x2[9] ),
    .S(net1952),
    .X(_00919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12749_ (.A0(\fpmul.reg_b_out[8] ),
    .A1(\fp16_res_pipe.x2[8] ),
    .S(net1955),
    .X(_00918_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12750_ (.A0(\fpmul.reg_b_out[7] ),
    .A1(\fp16_res_pipe.x2[7] ),
    .S(net1955),
    .X(_00917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12751_ (.Y(_06543_),
    .A(\fp16_res_pipe.x2[6] ),
    .B(net1955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12752_ (.B1(_06543_),
    .VDD(VPWR),
    .Y(_00916_),
    .VSS(VGND),
    .A1(net1956),
    .A2(_06031_));
 sg13g2_mux2_1 _12753_ (.A0(net1864),
    .A1(\fp16_res_pipe.x2[5] ),
    .S(net1957),
    .X(_00915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12754_ (.Y(_06544_),
    .A(\fp16_res_pipe.x2[4] ),
    .B(net1956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12755_ (.B1(_06544_),
    .VDD(VPWR),
    .Y(_00914_),
    .VSS(VGND),
    .A1(net1956),
    .A2(_06025_));
 sg13g2_mux2_1 _12756_ (.A0(\fpmul.reg_b_out[3] ),
    .A1(\fp16_res_pipe.x2[3] ),
    .S(net1957),
    .X(_00913_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12757_ (.Y(_06545_),
    .A(\fp16_res_pipe.x2[2] ),
    .B(net1957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12758_ (.B1(_06545_),
    .VDD(VPWR),
    .Y(_00912_),
    .VSS(VGND),
    .A1(net1957),
    .A2(_06015_));
 sg13g2_mux2_1 _12759_ (.A0(\fpmul.reg_b_out[1] ),
    .A1(\fp16_res_pipe.x2[1] ),
    .S(net1957),
    .X(_00911_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12760_ (.A0(\fpmul.reg_b_out[0] ),
    .A1(\fp16_res_pipe.x2[0] ),
    .S(net1957),
    .X(_00910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12761_ (.VDD(VPWR),
    .Y(_06546_),
    .A(net1941),
    .VSS(VGND));
 sg13g2_and3_1 _12762_ (.X(_06547_),
    .A(net1767),
    .B(\acc[15] ),
    .C(net1908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12763_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1909),
    .A2(\fp16_res_pipe.y[15] ),
    .Y(_06548_),
    .B1(_06547_));
 sg13g2_a21oi_1 _12764_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1923),
    .A2(\add_result[15] ),
    .Y(_06549_),
    .B1(net1941));
 sg13g2_o21ai_1 _12765_ (.B1(_06549_),
    .VDD(VPWR),
    .Y(_06550_),
    .VSS(VGND),
    .A1(net1923),
    .A2(_06548_));
 sg13g2_o21ai_1 _12766_ (.B1(_06550_),
    .VDD(VPWR),
    .Y(_06551_),
    .VSS(VGND),
    .A1(_06546_),
    .A2(\div_result[15] ));
 sg13g2_nor4_1 _12767_ (.A(_00016_),
    .B(_00015_),
    .C(_00014_),
    .D(_00013_),
    .Y(_06552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _12768_ (.A(_00020_),
    .B(_00019_),
    .C(_00018_),
    .D(_00017_),
    .Y(_06553_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _12769_ (.A(_00008_),
    .B(_00007_),
    .C(_00006_),
    .D(_00005_),
    .Y(_06554_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _12770_ (.A(_00012_),
    .B(_00011_),
    .C(_00010_),
    .D(_00009_),
    .Y(_06555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _12771_ (.B(_06553_),
    .C(_06554_),
    .A(_06552_),
    .Y(_06556_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_06555_));
 sg13g2_nor4_1 _12772_ (.A(\fpmul.reg3en.q[0] ),
    .B(\fpdiv.reg2en.q[0] ),
    .C(\fp16_sum_pipe.reg4en.q[0] ),
    .D(load_en),
    .Y(_06557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12773_ (.Y(_06558_),
    .A(_06557_),
    .B(_02623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _12774_ (.A(_06556_),
    .B_N(_06558_),
    .Y(_06559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout91 (.A(net92),
    .X(net91),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _12776_ (.Y(_06561_),
    .A(_06559_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12777_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1958),
    .A2(\fpmul.reg_p_out[15] ),
    .Y(_06562_),
    .B1(_06561_));
 sg13g2_o21ai_1 _12778_ (.B1(_06562_),
    .VDD(VPWR),
    .Y(_06563_),
    .VSS(VGND),
    .A1(net1958),
    .A2(_06551_));
 sg13g2_inv_1 _12779_ (.VDD(VPWR),
    .Y(_06564_),
    .A(\piso.tx_active ),
    .VSS(VGND));
 sg13g2_nor2_1 _12780_ (.A(net3),
    .B(_06564_),
    .Y(_06565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12781_ (.Y(_06566_),
    .A(_06561_),
    .B(_06565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12782_ (.VDD(VPWR),
    .Y(_06567_),
    .A(_06566_),
    .VSS(VGND));
 sg13g2_inv_1 _12783_ (.VDD(VPWR),
    .Y(_06568_),
    .A(\piso.tx_bit_counter[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12784_ (.Y(_06569_),
    .A(\piso.tx_bit_counter[1] ),
    .B(\piso.tx_bit_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12785_ (.A(_06568_),
    .B(_06569_),
    .Y(_06570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12786_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06570_),
    .A2(\piso.tx_bit_counter[3] ),
    .Y(_06571_),
    .B1(\piso.tx_bit_counter[4] ));
 sg13g2_buf_2 place1739 (.A(_02726_),
    .X(net1739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12788_ (.Y(_06573_),
    .A(_06567_),
    .B(_06571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _12789_ (.A(_06565_),
    .B(_06559_),
    .Y(_06574_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout110 (.A(net111),
    .X(net110),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout109 (.A(net113),
    .X(net109),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12792_ (.Y(_06577_),
    .A(net1716),
    .B(_00020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12793_ (.B(_06573_),
    .C(_06577_),
    .A(_06563_),
    .Y(_00909_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout127 (.A(net128),
    .X(net127),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1741 (.A(_02648_),
    .X(net1741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12796_ (.B(_00020_),
    .C(net1730),
    .A(net1701),
    .Y(_06580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12797_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[14] ),
    .Y(_06581_),
    .B1(net1943));
 sg13g2_nand3_1 _12798_ (.B(\acc[14] ),
    .C(net1908),
    .A(net1767),
    .Y(_06582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12799_ (.Y(_06583_),
    .A(net1910),
    .B(\fp16_res_pipe.y[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _12800_ (.A2(_06583_),
    .A1(_06582_),
    .B1(net1923),
    .X(_06584_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12801_ (.Y(_06585_),
    .B1(_06581_),
    .B2(_06584_),
    .A2(_06371_),
    .A1(net1941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12802_ (.VDD(VPWR),
    .Y(_06586_),
    .A(\fpmul.reg_p_out[14] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12803_ (.Y(_06587_),
    .A(_06586_),
    .B(net1958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12804_ (.B1(_06587_),
    .VDD(VPWR),
    .Y(_06588_),
    .VSS(VGND),
    .A1(net1958),
    .A2(_06585_));
 sg13g2_buf_2 fanout90 (.A(net91),
    .X(net90),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12806_ (.Y(_06590_),
    .A(_06588_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12807_ (.Y(_06591_),
    .A(net1716),
    .B(_00019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12808_ (.B(_06590_),
    .C(_06591_),
    .A(_06580_),
    .Y(_00908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12809_ (.B(_00019_),
    .C(net1730),
    .A(net1701),
    .Y(_06592_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12810_ (.VDD(VPWR),
    .Y(_06593_),
    .A(\div_result[13] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _12811_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[13] ),
    .Y(_06594_),
    .B1(net1943));
 sg13g2_nand3_1 _12812_ (.B(\acc[13] ),
    .C(net1908),
    .A(net1767),
    .Y(_06595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12813_ (.Y(_06596_),
    .A(net1909),
    .B(\fp16_res_pipe.y[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _12814_ (.A2(_06596_),
    .A1(_06595_),
    .B1(net1923),
    .X(_06597_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12815_ (.Y(_06598_),
    .B1(_06594_),
    .B2(_06597_),
    .A2(_06593_),
    .A1(net1941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12816_ (.VDD(VPWR),
    .Y(_06599_),
    .A(\fpmul.reg_p_out[13] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12817_ (.Y(_06600_),
    .A(_06599_),
    .B(net1959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12818_ (.B1(_06600_),
    .VDD(VPWR),
    .Y(_06601_),
    .VSS(VGND),
    .A1(net1960),
    .A2(_06598_));
 sg13g2_nand2_1 _12819_ (.Y(_06602_),
    .A(_06601_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12820_ (.Y(_06603_),
    .A(net1716),
    .B(_00018_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12821_ (.B(_06602_),
    .C(_06603_),
    .A(_06592_),
    .Y(_00907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12822_ (.B(_00018_),
    .C(net1730),
    .A(net1701),
    .Y(_06604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12823_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[12] ),
    .Y(_06605_),
    .B1(net1943));
 sg13g2_a21oi_1 _12824_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc[12] ),
    .A2(net1908),
    .Y(_06606_),
    .B1(net1909));
 sg13g2_a21oi_1 _12825_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04902_),
    .A2(net1911),
    .Y(_06607_),
    .B1(net1924));
 sg13g2_nand2b_1 _12826_ (.Y(_06608_),
    .B(_06607_),
    .A_N(_06606_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12827_ (.Y(_06609_),
    .B1(_06605_),
    .B2(_06608_),
    .A2(_06485_),
    .A1(net1941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12828_ (.VDD(VPWR),
    .Y(_06610_),
    .A(\fpmul.reg_p_out[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12829_ (.Y(_06611_),
    .A(_06610_),
    .B(net1959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12830_ (.B1(_06611_),
    .VDD(VPWR),
    .Y(_06612_),
    .VSS(VGND),
    .A1(net1958),
    .A2(_06609_));
 sg13g2_nand2_1 _12831_ (.Y(_06613_),
    .A(_06612_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12832_ (.Y(_06614_),
    .A(net1716),
    .B(_00017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12833_ (.B(_06613_),
    .C(_06614_),
    .A(_06604_),
    .Y(_00906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12834_ (.B(_00017_),
    .C(net1730),
    .A(net1701),
    .Y(_06615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12835_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[11] ),
    .Y(_06616_),
    .B1(net1943));
 sg13g2_nand3_1 _12836_ (.B(\acc[11] ),
    .C(net1908),
    .A(net1767),
    .Y(_06617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12837_ (.Y(_06618_),
    .A(net1909),
    .B(\fp16_res_pipe.y[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12838_ (.A2(_06618_),
    .A1(_06617_),
    .B1(net1922),
    .X(_06619_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12839_ (.Y(_06620_),
    .B1(_06616_),
    .B2(_06619_),
    .A2(_06488_),
    .A1(net1941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12840_ (.VDD(VPWR),
    .Y(_06621_),
    .A(\fpmul.reg_p_out[11] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12841_ (.Y(_06622_),
    .A(_06621_),
    .B(net1960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12842_ (.B1(_06622_),
    .VDD(VPWR),
    .Y(_06623_),
    .VSS(VGND),
    .A1(net1960),
    .A2(_06620_));
 sg13g2_nand2_1 _12843_ (.Y(_06624_),
    .A(_06623_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12844_ (.Y(_06625_),
    .A(net1716),
    .B(_00016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12845_ (.B(_06624_),
    .C(_06625_),
    .A(_06615_),
    .Y(_00905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12846_ (.B(_00016_),
    .C(net1730),
    .A(net1701),
    .Y(_06626_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12847_ (.VDD(VPWR),
    .Y(_06627_),
    .A(\div_result[10] ),
    .VSS(VGND));
 sg13g2_a21oi_1 _12848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[10] ),
    .Y(_06628_),
    .B1(net1943));
 sg13g2_a21oi_1 _12849_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc[10] ),
    .A2(net1907),
    .Y(_06629_),
    .B1(\fp16_res_pipe.reg1en.d[0] ));
 sg13g2_a21oi_1 _12850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04929_),
    .A2(net1911),
    .Y(_06630_),
    .B1(net1924));
 sg13g2_nand2b_1 _12851_ (.Y(_06631_),
    .B(_06630_),
    .A_N(_06629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12852_ (.Y(_06632_),
    .B1(_06628_),
    .B2(_06631_),
    .A2(_06627_),
    .A1(net1943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12853_ (.VDD(VPWR),
    .Y(_06633_),
    .A(\fpmul.reg_p_out[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12854_ (.Y(_06634_),
    .A(_06633_),
    .B(net1960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12855_ (.B1(_06634_),
    .VDD(VPWR),
    .Y(_06635_),
    .VSS(VGND),
    .A1(net1960),
    .A2(_06632_));
 sg13g2_nand2_1 _12856_ (.Y(_06636_),
    .A(_06635_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12857_ (.Y(_06637_),
    .A(_06574_),
    .B(_00015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12858_ (.B(_06636_),
    .C(_06637_),
    .A(_06626_),
    .Y(_00904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12859_ (.B(_00015_),
    .C(net1730),
    .A(net1701),
    .Y(_06638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[9] ),
    .Y(_06639_),
    .B1(net1943));
 sg13g2_a21oi_1 _12861_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\acc[9] ),
    .A2(net1907),
    .Y(_06640_),
    .B1(net1909));
 sg13g2_a21oi_1 _12862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_04940_),
    .A2(net1910),
    .Y(_06641_),
    .B1(net1923));
 sg13g2_nand2b_2 _12863_ (.Y(_06642_),
    .B(_06641_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06640_));
 sg13g2_a22oi_1 _12864_ (.Y(_06643_),
    .B1(_06639_),
    .B2(_06642_),
    .A2(_06496_),
    .A1(net1943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12865_ (.VDD(VPWR),
    .Y(_06644_),
    .A(\fpmul.reg_p_out[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12866_ (.Y(_06645_),
    .A(_06644_),
    .B(\fpmul.reg1en.d[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12867_ (.B1(_06645_),
    .VDD(VPWR),
    .Y(_06646_),
    .VSS(VGND),
    .A1(net1960),
    .A2(_06643_));
 sg13g2_nand2_1 _12868_ (.Y(_06647_),
    .A(_06646_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12869_ (.Y(_06648_),
    .A(_06574_),
    .B(_00014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12870_ (.B(_06647_),
    .C(_06648_),
    .A(_06638_),
    .Y(_00903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12871_ (.B(_00014_),
    .C(net1730),
    .A(net1701),
    .Y(_06649_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12872_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1935),
    .A2(\add_result[8] ),
    .Y(_06650_),
    .B1(net1949));
 sg13g2_nand3_1 _12873_ (.B(\acc[8] ),
    .C(net1908),
    .A(net1767),
    .Y(_06651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12874_ (.Y(_06652_),
    .A(net1909),
    .B(\fp16_res_pipe.y[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12875_ (.A2(_06652_),
    .A1(_06651_),
    .B1(net1922),
    .X(_06653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12876_ (.Y(_06654_),
    .B1(_06650_),
    .B2(_06653_),
    .A2(_06499_),
    .A1(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12877_ (.VDD(VPWR),
    .Y(_06655_),
    .A(\fpmul.reg_p_out[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12878_ (.Y(_06656_),
    .A(_06655_),
    .B(\fpmul.reg1en.d[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12879_ (.B1(_06656_),
    .VDD(VPWR),
    .Y(_06657_),
    .VSS(VGND),
    .A1(\fpmul.reg1en.d[0] ),
    .A2(_06654_));
 sg13g2_nand2_1 _12880_ (.Y(_06658_),
    .A(_06657_),
    .B(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12881_ (.Y(_06659_),
    .A(_06574_),
    .B(_00013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12882_ (.B(_06658_),
    .C(_06659_),
    .A(_06649_),
    .Y(_00902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12883_ (.B(_00013_),
    .C(net1731),
    .A(net1702),
    .Y(_06660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[7] ),
    .Y(_06661_),
    .B1(net1950));
 sg13g2_nand3_1 _12885_ (.B(\acc[7] ),
    .C(net1907),
    .A(net1767),
    .Y(_06662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12886_ (.Y(_06663_),
    .A(net1909),
    .B(\fp16_res_pipe.y[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12887_ (.A2(_06663_),
    .A1(_06662_),
    .B1(net1922),
    .X(_06664_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12888_ (.Y(_06665_),
    .B1(_06661_),
    .B2(_06664_),
    .A2(_06502_),
    .A1(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12889_ (.VDD(VPWR),
    .Y(_06666_),
    .A(\fpmul.reg_p_out[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12890_ (.Y(_06667_),
    .A(_06666_),
    .B(\fpmul.reg1en.d[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12891_ (.B1(_06667_),
    .VDD(VPWR),
    .Y(_06668_),
    .VSS(VGND),
    .A1(net1962),
    .A2(_06665_));
 sg13g2_nand2_1 _12892_ (.Y(_06669_),
    .A(_06668_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12893_ (.Y(_06670_),
    .A(net1717),
    .B(_00012_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12894_ (.B(_06669_),
    .C(_06670_),
    .A(_06660_),
    .Y(_00901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12895_ (.B(_00012_),
    .C(net1731),
    .A(net1702),
    .Y(_06671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12896_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[6] ),
    .Y(_06672_),
    .B1(net1950));
 sg13g2_nand3_1 _12897_ (.B(\acc[6] ),
    .C(net1907),
    .A(_03983_),
    .Y(_06673_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12898_ (.Y(_06674_),
    .A(net1910),
    .B(\fp16_res_pipe.y[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12899_ (.A2(_06674_),
    .A1(_06673_),
    .B1(\fp16_sum_pipe.reg1en.d[0] ),
    .X(_06675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12900_ (.Y(_06676_),
    .B1(_06672_),
    .B2(_06675_),
    .A2(_06510_),
    .A1(net1948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12901_ (.VDD(VPWR),
    .Y(_06677_),
    .A(\fpmul.reg_p_out[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12902_ (.Y(_06678_),
    .A(_06677_),
    .B(net1962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12903_ (.B1(_06678_),
    .VDD(VPWR),
    .Y(_06679_),
    .VSS(VGND),
    .A1(net1962),
    .A2(_06676_));
 sg13g2_nand2_1 _12904_ (.Y(_06680_),
    .A(_06679_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12905_ (.Y(_06681_),
    .A(net1717),
    .B(_00011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12906_ (.B(_06680_),
    .C(_06681_),
    .A(_06671_),
    .Y(_00900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12907_ (.B(_00011_),
    .C(net1731),
    .A(net1702),
    .Y(_06682_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[5] ),
    .Y(_06683_),
    .B1(net1950));
 sg13g2_nand3_1 _12909_ (.B(\acc[5] ),
    .C(net1908),
    .A(net1767),
    .Y(_06684_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12910_ (.Y(_06685_),
    .A(net1909),
    .B(\fp16_res_pipe.y[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12911_ (.A2(_06685_),
    .A1(_06684_),
    .B1(net1922),
    .X(_06686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12912_ (.Y(_06687_),
    .B1(_06683_),
    .B2(_06686_),
    .A2(_06516_),
    .A1(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12913_ (.VDD(VPWR),
    .Y(_06688_),
    .A(\fpmul.reg_p_out[5] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12914_ (.Y(_06689_),
    .A(_06688_),
    .B(net1961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12915_ (.B1(_06689_),
    .VDD(VPWR),
    .Y(_06690_),
    .VSS(VGND),
    .A1(net1962),
    .A2(_06687_));
 sg13g2_nand2_1 _12916_ (.Y(_06691_),
    .A(_06690_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12917_ (.Y(_06692_),
    .A(net1717),
    .B(_00010_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12918_ (.B(_06691_),
    .C(_06692_),
    .A(_06682_),
    .Y(_00899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12919_ (.B(_00010_),
    .C(net1731),
    .A(net1702),
    .Y(_06693_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[4] ),
    .Y(_06694_),
    .B1(net1950));
 sg13g2_nand3_1 _12921_ (.B(\acc[4] ),
    .C(net1907),
    .A(_03983_),
    .Y(_06695_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12922_ (.Y(_06696_),
    .A(\fp16_res_pipe.reg1en.d[0] ),
    .B(\fp16_res_pipe.y[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12923_ (.A2(_06696_),
    .A1(_06695_),
    .B1(net1922),
    .X(_06697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12924_ (.Y(_06698_),
    .B1(_06694_),
    .B2(_06697_),
    .A2(_06520_),
    .A1(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12925_ (.VDD(VPWR),
    .Y(_06699_),
    .A(\fpmul.reg_p_out[4] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12926_ (.Y(_06700_),
    .A(_06699_),
    .B(net1961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12927_ (.B1(_06700_),
    .VDD(VPWR),
    .Y(_06701_),
    .VSS(VGND),
    .A1(net1962),
    .A2(_06698_));
 sg13g2_nand2_1 _12928_ (.Y(_06702_),
    .A(_06701_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12929_ (.Y(_06703_),
    .A(net1717),
    .B(_00009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12930_ (.B(_06702_),
    .C(_06703_),
    .A(_06693_),
    .Y(_00898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12931_ (.B(_00009_),
    .C(net1731),
    .A(net1702),
    .Y(_06704_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12932_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[3] ),
    .Y(_06705_),
    .B1(net1950));
 sg13g2_nand3_1 _12933_ (.B(\acc[3] ),
    .C(net1907),
    .A(_03983_),
    .Y(_06706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12934_ (.Y(_06707_),
    .A(net1910),
    .B(\fp16_res_pipe.y[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12935_ (.A2(_06707_),
    .A1(_06706_),
    .B1(\fp16_sum_pipe.reg1en.d[0] ),
    .X(_06708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12936_ (.Y(_06709_),
    .B1(_06705_),
    .B2(_06708_),
    .A2(_06527_),
    .A1(net1948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12937_ (.VDD(VPWR),
    .Y(_06710_),
    .A(\fpmul.reg_p_out[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12938_ (.Y(_06711_),
    .A(_06710_),
    .B(net1962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12939_ (.B1(_06711_),
    .VDD(VPWR),
    .Y(_06712_),
    .VSS(VGND),
    .A1(net1962),
    .A2(_06709_));
 sg13g2_nand2_1 _12940_ (.Y(_06713_),
    .A(_06712_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12941_ (.Y(_06714_),
    .A(net1717),
    .B(_00008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12942_ (.B(_06713_),
    .C(_06714_),
    .A(_06704_),
    .Y(_00897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12943_ (.B(_00008_),
    .C(net1731),
    .A(net1702),
    .Y(_06715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[2] ),
    .Y(_06716_),
    .B1(net1950));
 sg13g2_nand3_1 _12945_ (.B(\acc[2] ),
    .C(load_en),
    .A(_03983_),
    .Y(_06717_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _12946_ (.Y(_06718_),
    .A(net1910),
    .B(\fp16_res_pipe.y[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12947_ (.A2(_06718_),
    .A1(_06717_),
    .B1(\fp16_sum_pipe.reg1en.d[0] ),
    .X(_06719_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12948_ (.Y(_06720_),
    .B1(_06716_),
    .B2(_06719_),
    .A2(_06533_),
    .A1(net1948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12949_ (.VDD(VPWR),
    .Y(_06721_),
    .A(\fpmul.reg_p_out[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12950_ (.Y(_06722_),
    .A(_06721_),
    .B(net1961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12951_ (.B1(_06722_),
    .VDD(VPWR),
    .Y(_06723_),
    .VSS(VGND),
    .A1(net1961),
    .A2(_06720_));
 sg13g2_nand2_1 _12952_ (.Y(_06724_),
    .A(_06723_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12953_ (.Y(_06725_),
    .A(net1717),
    .B(_00007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12954_ (.B(_06724_),
    .C(_06725_),
    .A(_06715_),
    .Y(_00896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12955_ (.B(_00007_),
    .C(net1731),
    .A(net1702),
    .Y(_06726_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[1] ),
    .Y(_06727_),
    .B1(net1950));
 sg13g2_nand3_1 _12957_ (.B(\acc[1] ),
    .C(load_en),
    .A(_03983_),
    .Y(_06728_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12958_ (.Y(_06729_),
    .A(net1910),
    .B(\fp16_res_pipe.y[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12959_ (.A2(_06729_),
    .A1(_06728_),
    .B1(\fp16_sum_pipe.reg1en.d[0] ),
    .X(_06730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12960_ (.Y(_06731_),
    .B1(_06727_),
    .B2(_06730_),
    .A2(_06536_),
    .A1(net1948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12961_ (.VDD(VPWR),
    .Y(_06732_),
    .A(\fpmul.reg_p_out[1] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12962_ (.Y(_06733_),
    .A(_06732_),
    .B(net1961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12963_ (.B1(_06733_),
    .VDD(VPWR),
    .Y(_06734_),
    .VSS(VGND),
    .A1(net1961),
    .A2(_06731_));
 sg13g2_nand2_1 _12964_ (.Y(_06735_),
    .A(_06734_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12965_ (.Y(_06736_),
    .A(net1717),
    .B(_00006_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12966_ (.B(_06735_),
    .C(_06736_),
    .A(_06726_),
    .Y(_00895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12967_ (.B(_00006_),
    .C(net1731),
    .A(net1702),
    .Y(_06737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _12968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1936),
    .A2(\add_result[0] ),
    .Y(_06738_),
    .B1(net1950));
 sg13g2_nand3_1 _12969_ (.B(\acc[0] ),
    .C(net1907),
    .A(_03983_),
    .Y(_06739_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12970_ (.Y(_06740_),
    .A(net1910),
    .B(\fp16_res_pipe.y[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_2 _12971_ (.A2(_06740_),
    .A1(_06739_),
    .B1(\fp16_sum_pipe.reg1en.d[0] ),
    .X(_06741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _12972_ (.Y(_06742_),
    .B1(_06738_),
    .B2(_06741_),
    .A2(_06539_),
    .A1(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12973_ (.VDD(VPWR),
    .Y(_06743_),
    .A(\fpmul.reg_p_out[0] ),
    .VSS(VGND));
 sg13g2_nand2_1 _12974_ (.Y(_06744_),
    .A(_06743_),
    .B(net1961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _12975_ (.B1(_06744_),
    .VDD(VPWR),
    .Y(_06745_),
    .VSS(VGND),
    .A1(net1962),
    .A2(_06742_));
 sg13g2_nand2_1 _12976_ (.Y(_06746_),
    .A(_06745_),
    .B(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12977_ (.Y(_06747_),
    .A(net1717),
    .B(_00005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _12978_ (.B(_06746_),
    .C(_06747_),
    .A(_06737_),
    .Y(_00894_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _12979_ (.A0(\fpmul.reg_p_out[15] ),
    .A1(\fpmul.result[15] ),
    .S(net1861),
    .X(_00893_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12980_ (.VDD(VPWR),
    .Y(_06748_),
    .A(\fpmul.seg_reg0.q[22] ),
    .VSS(VGND));
 sg13g2_inv_1 _12981_ (.VDD(VPWR),
    .Y(_06749_),
    .A(\fpmul.seg_reg0.q[20] ),
    .VSS(VGND));
 sg13g2_inv_2 _12982_ (.Y(_06750_),
    .A(\fpmul.seg_reg0.q[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _12983_ (.A(_05873_),
    .B(_05877_),
    .C(net1755),
    .Y(_06751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _12984_ (.Y(_06752_),
    .A(_06751_),
    .B(\fpmul.seg_reg0.q[18] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _12985_ (.A(_05868_),
    .B(_06752_),
    .Y(_06753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12986_ (.VDD(VPWR),
    .Y(_06754_),
    .A(_06753_),
    .VSS(VGND));
 sg13g2_nor2_1 _12987_ (.A(_06749_),
    .B(_06754_),
    .Y(_06755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _12988_ (.Y(_06756_),
    .A(_05863_),
    .B(_06755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12989_ (.VDD(VPWR),
    .Y(_06757_),
    .A(_06756_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12990_ (.Y(_06758_),
    .A(_06749_),
    .B(_06753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12991_ (.VDD(VPWR),
    .Y(_06759_),
    .A(_06758_),
    .VSS(VGND));
 sg13g2_xnor2_1 _12992_ (.Y(_06760_),
    .A(\fpmul.seg_reg0.q[19] ),
    .B(_06752_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12993_ (.VDD(VPWR),
    .Y(_06761_),
    .A(_06760_),
    .VSS(VGND));
 sg13g2_xor2_1 _12994_ (.B(_06751_),
    .A(\fpmul.seg_reg0.q[18] ),
    .X(_06762_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12995_ (.VDD(VPWR),
    .Y(_06763_),
    .A(_06762_),
    .VSS(VGND));
 sg13g2_xor2_1 _12996_ (.B(\fpmul.seg_reg0.q[15] ),
    .A(\fpmul.seg_reg0.q[16] ),
    .X(_06764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _12997_ (.VDD(VPWR),
    .Y(_06765_),
    .A(_06764_),
    .VSS(VGND));
 sg13g2_nor2_1 _12998_ (.A(\fpmul.seg_reg0.q[15] ),
    .B(\fpmul.seg_reg0.q[14] ),
    .Y(_06766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _12999_ (.Y(_06767_),
    .B(net1755),
    .A_N(\fpmul.seg_reg0.q[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13000_ (.B1(_06767_),
    .VDD(VPWR),
    .Y(_06768_),
    .VSS(VGND),
    .A1(net1755),
    .A2(\fpmul.seg_reg0.q[14] ));
 sg13g2_nand2_1 _13001_ (.Y(_06769_),
    .A(\fpmul.seg_reg0.q[15] ),
    .B(\fpmul.seg_reg0.q[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13002_ (.VDD(VPWR),
    .Y(_06770_),
    .A(_06769_),
    .VSS(VGND));
 sg13g2_a21oi_1 _13003_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1755),
    .A2(\fpmul.seg_reg0.q[12] ),
    .Y(_06771_),
    .B1(_06770_));
 sg13g2_nand2_1 _13004_ (.Y(_06772_),
    .A(\fpmul.seg_reg0.q[15] ),
    .B(\fpmul.seg_reg0.q[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13005_ (.VDD(VPWR),
    .Y(_06773_),
    .A(_06772_),
    .VSS(VGND));
 sg13g2_a21oi_2 _13006_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_06773_),
    .Y(_06774_),
    .A2(\fpmul.seg_reg0.q[11] ),
    .A1(net1755));
 sg13g2_nor2_1 _13007_ (.A(net1853),
    .B(\fpmul.seg_reg0.q[7] ),
    .Y(_06775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _13008_ (.Y(_06776_),
    .B(net1853),
    .A_N(\fpmul.seg_reg0.q[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _13009_ (.Y(_06777_),
    .B(_06776_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06775_));
 sg13g2_nand2b_1 _13010_ (.Y(_06778_),
    .B(_06750_),
    .A_N(\fpmul.seg_reg0.q[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13011_ (.B1(_06778_),
    .VDD(VPWR),
    .Y(_06779_),
    .VSS(VGND),
    .A1(_06750_),
    .A2(\fpmul.seg_reg0.q[9] ));
 sg13g2_buf_2 place1738 (.A(_03365_),
    .X(net1738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13013_ (.A(_06777_),
    .B(_06779_),
    .Y(_06781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13014_ (.A(net1853),
    .B(\fpmul.seg_reg0.q[9] ),
    .Y(_06782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _13015_ (.A2(_06313_),
    .A1(net1853),
    .B1(_06782_),
    .X(_06783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13016_ (.VDD(VPWR),
    .Y(_06784_),
    .A(_06783_),
    .VSS(VGND));
 sg13g2_nand2_1 _13017_ (.Y(_06785_),
    .A(_06304_),
    .B(net1853),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13018_ (.B1(_06785_),
    .VDD(VPWR),
    .Y(_06786_),
    .VSS(VGND),
    .A1(net1853),
    .A2(\fpmul.seg_reg0.q[10] ));
 sg13g2_inv_1 _13019_ (.VDD(VPWR),
    .Y(_06787_),
    .A(_06786_),
    .VSS(VGND));
 sg13g2_nand3_1 _13020_ (.B(_06784_),
    .C(_06787_),
    .A(_06781_),
    .Y(_06788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout120 (.A(net122),
    .X(net120),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _13022_ (.A(_06771_),
    .B(_06774_),
    .C(_06788_),
    .Y(_06790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13023_ (.VDD(VPWR),
    .Y(_06791_),
    .A(_06790_),
    .VSS(VGND));
 sg13g2_nor3_1 _13024_ (.A(_06766_),
    .B(_06768_),
    .C(_06791_),
    .Y(_06792_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13025_ (.Y(_06793_),
    .A(net1853),
    .B(\fpmul.seg_reg0.q[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13026_ (.VDD(VPWR),
    .Y(_06794_),
    .A(_06793_),
    .VSS(VGND));
 sg13g2_a21oi_1 _13027_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1755),
    .A2(\fpmul.seg_reg0.q[6] ),
    .Y(_06795_),
    .B1(_06794_));
 sg13g2_inv_1 _13028_ (.VDD(VPWR),
    .Y(_06796_),
    .A(_06795_),
    .VSS(VGND));
 sg13g2_nand2_1 _13029_ (.Y(_06797_),
    .A(net1853),
    .B(\fpmul.seg_reg0.q[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13030_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06750_),
    .A2(\fpmul.seg_reg0.q[4] ),
    .Y(_06798_),
    .B1(\fpmul.seg_reg0.q[5] ));
 sg13g2_and3_1 _13031_ (.X(_06799_),
    .A(_06796_),
    .B(_06797_),
    .C(_06798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _13032_ (.A(_06799_),
    .B(_06777_),
    .X(_06800_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _13033_ (.A(_06795_),
    .B(_06800_),
    .Y(_06801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _13034_ (.Y(_06802_),
    .A(_06792_),
    .B(_06801_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1684 (.A(_02250_),
    .X(net1684),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13036_ (.A(_06765_),
    .B(_06802_),
    .Y(_06804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13037_ (.VDD(VPWR),
    .Y(_06805_),
    .A(_06804_),
    .VSS(VGND));
 sg13g2_nor2_1 _13038_ (.A(_05873_),
    .B(_06805_),
    .Y(_06806_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13039_ (.VDD(VPWR),
    .Y(_06807_),
    .A(_06806_),
    .VSS(VGND));
 sg13g2_nor2_1 _13040_ (.A(_06763_),
    .B(_06807_),
    .Y(_06808_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13041_ (.VDD(VPWR),
    .Y(_06809_),
    .A(_06808_),
    .VSS(VGND));
 sg13g2_nor2_1 _13042_ (.A(_06761_),
    .B(_06809_),
    .Y(_06810_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13043_ (.VDD(VPWR),
    .Y(_06811_),
    .A(_06810_),
    .VSS(VGND));
 sg13g2_nor2_1 _13044_ (.A(_06759_),
    .B(_06811_),
    .Y(_06812_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13045_ (.VDD(VPWR),
    .Y(_06813_),
    .A(_06812_),
    .VSS(VGND));
 sg13g2_nor2_1 _13046_ (.A(_06757_),
    .B(_06813_),
    .Y(_06814_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13047_ (.VDD(VPWR),
    .Y(_06815_),
    .A(_06814_),
    .VSS(VGND));
 sg13g2_nor2_1 _13048_ (.A(_06748_),
    .B(_06815_),
    .Y(_06816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13049_ (.VDD(VPWR),
    .Y(_06817_),
    .A(_06816_),
    .VSS(VGND));
 sg13g2_nor3_1 _13050_ (.A(_05863_),
    .B(_06749_),
    .C(_06754_),
    .Y(_06818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13051_ (.Y(_06819_),
    .A(_06818_),
    .B(\fpmul.seg_reg0.q[22] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _13052_ (.B(_06819_),
    .A(\fpmul.seg_reg0.q[23] ),
    .X(_06820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13053_ (.Y(_06821_),
    .A(_06817_),
    .B(_06820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _13054_ (.A(\fpmul.seg_reg0.q[49] ),
    .B(\fpmul.seg_reg0.q[48] ),
    .C(\fpmul.seg_reg0.q[47] ),
    .D(\fpmul.seg_reg0.q[46] ),
    .Y(_06822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _13055_ (.A(\fpmul.seg_reg0.q[53] ),
    .B(\fpmul.seg_reg0.q[52] ),
    .C(\fpmul.seg_reg0.q[51] ),
    .Y(_06823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13056_ (.Y(_06824_),
    .A(_06822_),
    .B(_06823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _13057_ (.A(\fpmul.seg_reg0.q[45] ),
    .B(\fpmul.seg_reg0.q[44] ),
    .C(\fpmul.seg_reg0.q[43] ),
    .D(\fpmul.seg_reg0.q[42] ),
    .Y(_06825_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _13058_ (.B(_05787_),
    .C(_05789_),
    .A(_06825_),
    .Y(_06826_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05791_));
 sg13g2_nor3_1 _13059_ (.A(\fpmul.seg_reg0.q[50] ),
    .B(_06824_),
    .C(_06826_),
    .Y(_06827_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13060_ (.VDD(VPWR),
    .Y(_06828_),
    .A(_06827_),
    .VSS(VGND));
 sg13g2_nand3_1 _13061_ (.B(_05813_),
    .C(_05819_),
    .A(_05811_),
    .Y(_06829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _13062_ (.B(_05803_),
    .C(_05805_),
    .A(_05801_),
    .Y(_06830_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05807_));
 sg13g2_nand4_1 _13063_ (.B(_05795_),
    .C(_05797_),
    .A(_05793_),
    .Y(_06831_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05799_));
 sg13g2_nand4_1 _13064_ (.B(_05815_),
    .C(_05817_),
    .A(_05809_),
    .Y(_06832_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_05821_));
 sg13g2_nor4_1 _13065_ (.A(_06829_),
    .B(_06830_),
    .C(_06831_),
    .D(_06832_),
    .Y(_06833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13066_ (.VDD(VPWR),
    .Y(_06834_),
    .A(_06833_),
    .VSS(VGND));
 sg13g2_nand3_1 _13067_ (.B(\fpmul.reg2en.q[0] ),
    .C(_06834_),
    .A(_06828_),
    .Y(_06835_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1751 (.A(_06903_),
    .X(net1751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13069_ (.VDD(VPWR),
    .Y(_06837_),
    .A(_06835_),
    .VSS(VGND));
 sg13g2_nand2b_1 _13070_ (.Y(_06838_),
    .B(_06816_),
    .A_N(_06820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13071_ (.B(_06837_),
    .C(_06838_),
    .A(_06821_),
    .Y(_06839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13072_ (.B1(_06839_),
    .VDD(VPWR),
    .Y(_00892_),
    .VSS(VGND),
    .A1(net1861),
    .A2(_06586_));
 sg13g2_nand2b_1 _13073_ (.Y(_06840_),
    .B(_06748_),
    .A_N(_06818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13074_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06819_),
    .A2(_06840_),
    .Y(_06841_),
    .B1(_06814_));
 sg13g2_nand3b_1 _13075_ (.B(_06817_),
    .C(_06837_),
    .Y(_06842_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06841_));
 sg13g2_o21ai_1 _13076_ (.B1(_06842_),
    .VDD(VPWR),
    .Y(_00891_),
    .VSS(VGND),
    .A1(net1861),
    .A2(_06599_));
 sg13g2_a21oi_1 _13077_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06813_),
    .A2(_06757_),
    .Y(_06843_),
    .B1(_06835_));
 sg13g2_nand2_1 _13078_ (.Y(_06844_),
    .A(_06843_),
    .B(_06815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13079_ (.B1(_06844_),
    .VDD(VPWR),
    .Y(_00890_),
    .VSS(VGND),
    .A1(net1861),
    .A2(_06610_));
 sg13g2_a21oi_1 _13080_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06811_),
    .A2(_06759_),
    .Y(_06845_),
    .B1(_06835_));
 sg13g2_nand2_1 _13081_ (.Y(_06846_),
    .A(_06845_),
    .B(_06813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13082_ (.B1(_06846_),
    .VDD(VPWR),
    .Y(_00889_),
    .VSS(VGND),
    .A1(net1861),
    .A2(_06621_));
 sg13g2_a21oi_1 _13083_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06809_),
    .A2(_06761_),
    .Y(_06847_),
    .B1(_06835_));
 sg13g2_nand2_1 _13084_ (.Y(_06848_),
    .A(_06847_),
    .B(_06811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13085_ (.B1(_06848_),
    .VDD(VPWR),
    .Y(_00888_),
    .VSS(VGND),
    .A1(net1861),
    .A2(_06633_));
 sg13g2_nand2_1 _13086_ (.Y(_06849_),
    .A(_06807_),
    .B(_06763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13087_ (.B(net1700),
    .C(_06849_),
    .A(_06809_),
    .Y(_06850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13088_ (.B1(_06850_),
    .VDD(VPWR),
    .Y(_00887_),
    .VSS(VGND),
    .A1(net1861),
    .A2(_06644_));
 sg13g2_a21oi_1 _13089_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\fpmul.seg_reg0.q[16] ),
    .A2(\fpmul.seg_reg0.q[15] ),
    .Y(_06851_),
    .B1(\fpmul.seg_reg0.q[17] ));
 sg13g2_o21ai_1 _13090_ (.B1(_06805_),
    .VDD(VPWR),
    .Y(_06852_),
    .VSS(VGND),
    .A1(_06751_),
    .A2(_06851_));
 sg13g2_nand3_1 _13091_ (.B(_06807_),
    .C(net1700),
    .A(_06852_),
    .Y(_06853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13092_ (.B1(_06853_),
    .VDD(VPWR),
    .Y(_00886_),
    .VSS(VGND),
    .A1(\fpmul.reg2en.q[0] ),
    .A2(_06655_));
 sg13g2_a21oi_1 _13093_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06802_),
    .A2(_06765_),
    .Y(_06854_),
    .B1(_06835_));
 sg13g2_nand2_1 _13094_ (.Y(_06855_),
    .A(_06854_),
    .B(_06805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13095_ (.B1(_06855_),
    .VDD(VPWR),
    .Y(_00885_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06666_));
 sg13g2_inv_1 _13096_ (.VDD(VPWR),
    .Y(_06856_),
    .A(_06801_),
    .VSS(VGND));
 sg13g2_o21ai_1 _13097_ (.B1(_06768_),
    .VDD(VPWR),
    .Y(_06857_),
    .VSS(VGND),
    .A1(_06791_),
    .A2(_06856_));
 sg13g2_nand3b_1 _13098_ (.B(_06801_),
    .C(_06790_),
    .Y(_06858_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06768_));
 sg13g2_nand3_1 _13099_ (.B(net1700),
    .C(_06858_),
    .A(_06857_),
    .Y(_06859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13100_ (.B1(_06859_),
    .VDD(VPWR),
    .Y(_00884_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06677_));
 sg13g2_o21ai_1 _13101_ (.B1(_06771_),
    .VDD(VPWR),
    .Y(_06860_),
    .VSS(VGND),
    .A1(_06774_),
    .A2(_06788_));
 sg13g2_nand3_1 _13102_ (.B(_06860_),
    .C(_06791_),
    .A(_06801_),
    .Y(_06861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13103_ (.B1(_06861_),
    .VDD(VPWR),
    .Y(_06862_),
    .VSS(VGND),
    .A1(_06771_),
    .A2(_06801_));
 sg13g2_nand3_1 _13104_ (.B(_06802_),
    .C(net1700),
    .A(_06862_),
    .Y(_06863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13105_ (.B1(_06863_),
    .VDD(VPWR),
    .Y(_00883_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06688_));
 sg13g2_a21oi_1 _13106_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06774_),
    .A2(_06856_),
    .Y(_06864_),
    .B1(_06835_));
 sg13g2_xor2_1 _13107_ (.B(_06788_),
    .A(_06774_),
    .X(_06865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _13108_ (.Y(_06866_),
    .B(_06801_),
    .A_N(_06865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13109_ (.B(_06802_),
    .C(_06866_),
    .A(_06864_),
    .Y(_06867_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13110_ (.B1(_06867_),
    .VDD(VPWR),
    .Y(_00882_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06699_));
 sg13g2_nand2b_2 _13111_ (.Y(_06868_),
    .B(_06796_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_06777_));
 sg13g2_nor2_1 _13112_ (.A(_06779_),
    .B(_06868_),
    .Y(_06869_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13113_ (.Y(_06870_),
    .A(_06869_),
    .B(_06784_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _13114_ (.Y(_06871_),
    .A(_06787_),
    .B(_06870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13115_ (.B(net1700),
    .C(_06871_),
    .A(_06802_),
    .Y(_06872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13116_ (.B1(_06872_),
    .VDD(VPWR),
    .Y(_00881_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06710_));
 sg13g2_o21ai_1 _13117_ (.B1(_06783_),
    .VDD(VPWR),
    .Y(_06873_),
    .VSS(VGND),
    .A1(_06779_),
    .A2(_06868_));
 sg13g2_nand4_1 _13118_ (.B(net1700),
    .C(_06870_),
    .A(_06802_),
    .Y(_06874_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_06873_));
 sg13g2_o21ai_1 _13119_ (.B1(_06874_),
    .VDD(VPWR),
    .Y(_00880_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06721_));
 sg13g2_xor2_1 _13120_ (.B(_06868_),
    .A(_06779_),
    .X(_06875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13121_ (.B(net1700),
    .C(_06875_),
    .A(_06802_),
    .Y(_06876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13122_ (.B1(_06876_),
    .VDD(VPWR),
    .Y(_00879_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06732_));
 sg13g2_or2_1 _13123_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_06877_),
    .B(_06792_),
    .A(_06868_));
 sg13g2_o21ai_1 _13124_ (.B1(_06777_),
    .VDD(VPWR),
    .Y(_06878_),
    .VSS(VGND),
    .A1(_06795_),
    .A2(_06799_));
 sg13g2_nand4_1 _13125_ (.B(_06802_),
    .C(net1700),
    .A(_06877_),
    .Y(_06879_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_06878_));
 sg13g2_o21ai_1 _13126_ (.B1(_06879_),
    .VDD(VPWR),
    .Y(_00878_),
    .VSS(VGND),
    .A1(net1862),
    .A2(_06743_));
 sg13g2_inv_4 _13127_ (.A(net3),
    .Y(_06880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13128_ (.B1(_06880_),
    .VDD(VPWR),
    .Y(_06881_),
    .VSS(VGND),
    .A1(_06564_),
    .A2(_06558_));
 sg13g2_or2_1 _13129_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_06882_),
    .B(_06881_),
    .A(_06556_));
 sg13g2_buf_2 place1735 (.A(net1734),
    .X(net1735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _13131_ (.A(_06882_),
    .B_N(\piso.tx_bit_counter[4] ),
    .Y(_00877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13132_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06882_),
    .A2(_06570_),
    .Y(_06884_),
    .B1(\piso.tx_bit_counter[3] ));
 sg13g2_nand2_1 _13133_ (.Y(_06885_),
    .A(_06573_),
    .B(_06882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13134_ (.VDD(VPWR),
    .Y(_06886_),
    .A(_06885_),
    .VSS(VGND));
 sg13g2_nor2_1 _13135_ (.A(_06884_),
    .B(_06886_),
    .Y(_00876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _13136_ (.A(_06569_),
    .B_N(_06882_),
    .Y(_06887_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13137_ (.VDD(VPWR),
    .Y(_06888_),
    .A(_06887_),
    .VSS(VGND));
 sg13g2_nand3_1 _13138_ (.B(_06564_),
    .C(_06880_),
    .A(_06556_),
    .Y(_06889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13139_ (.VDD(VPWR),
    .Y(_06890_),
    .A(_06889_),
    .VSS(VGND));
 sg13g2_nor3_1 _13140_ (.A(\piso.tx_bit_counter[4] ),
    .B(net3),
    .C(_06890_),
    .Y(_06891_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _13141_ (.Y(_06892_),
    .B(_06891_),
    .A_N(_06570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _13142_ (.Y(_00875_),
    .B1(_06882_),
    .B2(_06892_),
    .A2(_06888_),
    .A1(_06568_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13143_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06882_),
    .A2(\piso.tx_bit_counter[0] ),
    .Y(_06893_),
    .B1(\piso.tx_bit_counter[1] ));
 sg13g2_nor3_1 _13144_ (.A(_06887_),
    .B(_06893_),
    .C(_06886_),
    .Y(_00874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13145_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06891_),
    .A2(_06882_),
    .Y(_06894_),
    .B1(\piso.tx_bit_counter[0] ));
 sg13g2_a21oi_1 _13146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\piso.tx_bit_counter[0] ),
    .A2(_06882_),
    .Y(_00873_),
    .B1(_06894_));
 sg13g2_nand2_1 _13147_ (.Y(_06895_),
    .A(_06566_),
    .B(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13148_ (.B1(_06895_),
    .VDD(VPWR),
    .Y(_00872_),
    .VSS(VGND),
    .A1(_00005_),
    .A2(_06566_));
 sg13g2_nand2_1 _13149_ (.Y(_06896_),
    .A(_06885_),
    .B(\piso.tx_active ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13150_ (.Y(_00871_),
    .A(_06896_),
    .B(_06889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13151_ (.VDD(VPWR),
    .Y(_06897_),
    .A(\sipo.bit_counter[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13152_ (.Y(_06898_),
    .A(\sipo.bit_counter[1] ),
    .B(\sipo.bit_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13153_ (.A(_06897_),
    .B(_06898_),
    .Y(_06899_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13154_ (.Y(_06900_),
    .A(_06899_),
    .B(\sipo.bit_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _13155_ (.A(\sipo.bit_counter[4] ),
    .B(_06900_),
    .Y(_06901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _13156_ (.Y(_06902_),
    .A(_06901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _13157_ (.Y(_06903_),
    .A(_06880_),
    .B(\sipo.receiving ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout63 (.A(net67),
    .X(net63),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _13159_ (.Y(_06905_),
    .A(_06903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13160_ (.Y(_06906_),
    .A(_06905_),
    .B(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _13161_ (.Y(_06907_),
    .A(_06901_),
    .B(_06905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout116 (.A(net119),
    .X(net116),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout115 (.A(net116),
    .X(net115),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13164_ (.Y(_06910_),
    .A(net1713),
    .B(\sipo.word[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13165_ (.B1(_06910_),
    .VDD(VPWR),
    .Y(_00870_),
    .VSS(VGND),
    .A1(_06902_),
    .A2(_06906_));
 sg13g2_inv_1 _13166_ (.VDD(VPWR),
    .Y(_06911_),
    .A(\sipo.shift_reg[15] ),
    .VSS(VGND));
 sg13g2_buf_2 fanout114 (.A(net116),
    .X(net114),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13168_ (.Y(_06913_),
    .A(net1713),
    .B(\sipo.word[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13169_ (.B1(_06913_),
    .VDD(VPWR),
    .Y(_00869_),
    .VSS(VGND),
    .A1(_06911_),
    .A2(net1713));
 sg13g2_inv_1 _13170_ (.VDD(VPWR),
    .Y(_06914_),
    .A(\sipo.shift_reg[14] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13171_ (.Y(_06915_),
    .A(_06907_),
    .B(\sipo.word[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13172_ (.B1(_06915_),
    .VDD(VPWR),
    .Y(_00868_),
    .VSS(VGND),
    .A1(_06914_),
    .A2(_06907_));
 sg13g2_inv_1 _13173_ (.VDD(VPWR),
    .Y(_06916_),
    .A(\sipo.shift_reg[13] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13174_ (.Y(_06917_),
    .A(net1712),
    .B(\sipo.word[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13175_ (.B1(_06917_),
    .VDD(VPWR),
    .Y(_00867_),
    .VSS(VGND),
    .A1(_06916_),
    .A2(net1712));
 sg13g2_inv_1 _13176_ (.VDD(VPWR),
    .Y(_06918_),
    .A(\sipo.shift_reg[12] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13177_ (.Y(_06919_),
    .A(net1715),
    .B(\sipo.word[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13178_ (.B1(_06919_),
    .VDD(VPWR),
    .Y(_00866_),
    .VSS(VGND),
    .A1(_06918_),
    .A2(net1715));
 sg13g2_inv_1 _13179_ (.VDD(VPWR),
    .Y(_06920_),
    .A(\sipo.shift_reg[11] ),
    .VSS(VGND));
 sg13g2_buf_1 fanout113 (.A(net128),
    .X(net113),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13181_ (.Y(_06922_),
    .A(net1715),
    .B(\sipo.word[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13182_ (.B1(_06922_),
    .VDD(VPWR),
    .Y(_00865_),
    .VSS(VGND),
    .A1(_06920_),
    .A2(net1715));
 sg13g2_inv_1 _13183_ (.VDD(VPWR),
    .Y(_06923_),
    .A(\sipo.shift_reg[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13184_ (.Y(_06924_),
    .A(net1715),
    .B(\sipo.word[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13185_ (.B1(_06924_),
    .VDD(VPWR),
    .Y(_00864_),
    .VSS(VGND),
    .A1(_06923_),
    .A2(net1715));
 sg13g2_inv_1 _13186_ (.VDD(VPWR),
    .Y(_06925_),
    .A(\sipo.shift_reg[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13187_ (.Y(_06926_),
    .A(net1712),
    .B(\sipo.word[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13188_ (.B1(_06926_),
    .VDD(VPWR),
    .Y(_00863_),
    .VSS(VGND),
    .A1(_06925_),
    .A2(net1712));
 sg13g2_inv_1 _13189_ (.VDD(VPWR),
    .Y(_06927_),
    .A(\sipo.shift_reg[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13190_ (.Y(_06928_),
    .A(net1712),
    .B(\sipo.word[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13191_ (.B1(_06928_),
    .VDD(VPWR),
    .Y(_00862_),
    .VSS(VGND),
    .A1(_06927_),
    .A2(net1712));
 sg13g2_inv_1 _13192_ (.VDD(VPWR),
    .Y(_06929_),
    .A(\sipo.shift_reg[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13193_ (.Y(_06930_),
    .A(net1712),
    .B(\sipo.word[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13194_ (.B1(_06930_),
    .VDD(VPWR),
    .Y(_00861_),
    .VSS(VGND),
    .A1(_06929_),
    .A2(net1712));
 sg13g2_inv_1 _13195_ (.VDD(VPWR),
    .Y(_06931_),
    .A(\sipo.shift_reg[6] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13196_ (.Y(_06932_),
    .A(net1713),
    .B(\sipo.word[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13197_ (.B1(_06932_),
    .VDD(VPWR),
    .Y(_00860_),
    .VSS(VGND),
    .A1(_06931_),
    .A2(net1713));
 sg13g2_inv_1 _13198_ (.VDD(VPWR),
    .Y(_06933_),
    .A(\sipo.shift_reg[5] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13199_ (.Y(_06934_),
    .A(net1713),
    .B(\sipo.word[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13200_ (.B1(_06934_),
    .VDD(VPWR),
    .Y(_00859_),
    .VSS(VGND),
    .A1(_06933_),
    .A2(net1713));
 sg13g2_inv_1 _13201_ (.VDD(VPWR),
    .Y(_06935_),
    .A(\sipo.shift_reg[4] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13202_ (.Y(_06936_),
    .A(net1714),
    .B(\sipo.word[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13203_ (.B1(_06936_),
    .VDD(VPWR),
    .Y(_00858_),
    .VSS(VGND),
    .A1(_06935_),
    .A2(net1714));
 sg13g2_inv_1 _13204_ (.VDD(VPWR),
    .Y(_06937_),
    .A(\sipo.shift_reg[3] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13205_ (.Y(_06938_),
    .A(net1714),
    .B(\sipo.word[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13206_ (.B1(_06938_),
    .VDD(VPWR),
    .Y(_00857_),
    .VSS(VGND),
    .A1(_06937_),
    .A2(net1714));
 sg13g2_inv_1 _13207_ (.VDD(VPWR),
    .Y(_06939_),
    .A(\sipo.shift_reg[2] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13208_ (.Y(_06940_),
    .A(net1714),
    .B(\sipo.word[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13209_ (.B1(_06940_),
    .VDD(VPWR),
    .Y(_00856_),
    .VSS(VGND),
    .A1(_06939_),
    .A2(net1714));
 sg13g2_inv_2 _13210_ (.Y(_06941_),
    .A(\sipo.word[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13211_ (.A(\sipo.shift_reg[1] ),
    .B(net1714),
    .Y(_06942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13212_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06941_),
    .A2(net1714),
    .Y(_00855_),
    .B1(_06942_));
 sg13g2_a21oi_1 _13213_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06900_),
    .A2(\sipo.receiving ),
    .Y(_06943_),
    .B1(net3));
 sg13g2_nor2b_1 _13214_ (.A(_06943_),
    .B_N(\sipo.bit_counter[4] ),
    .Y(_00854_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13215_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06899_),
    .A2(_06880_),
    .Y(_06944_),
    .B1(\sipo.bit_counter[3] ));
 sg13g2_nor2_1 _13216_ (.A(_06944_),
    .B(_06943_),
    .Y(_00853_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13217_ (.VDD(VPWR),
    .Y(_06945_),
    .A(_06898_),
    .VSS(VGND));
 sg13g2_nor2_1 _13218_ (.A(_06903_),
    .B(_06899_),
    .Y(_06946_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13219_ (.B1(_06946_),
    .VDD(VPWR),
    .Y(_06947_),
    .VSS(VGND),
    .A1(\sipo.bit_counter[2] ),
    .A2(_06945_));
 sg13g2_o21ai_1 _13220_ (.B1(_06947_),
    .VDD(VPWR),
    .Y(_00852_),
    .VSS(VGND),
    .A1(_06897_),
    .A2(_06880_));
 sg13g2_nor2_1 _13221_ (.A(\sipo.bit_counter[1] ),
    .B(\sipo.bit_counter[0] ),
    .Y(_06948_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _13222_ (.A(_06948_),
    .B(_06903_),
    .C(_06945_),
    .Y(_06949_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _13223_ (.A2(net3),
    .A1(\sipo.bit_counter[1] ),
    .B1(_06949_),
    .X(_00851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout62 (.A(net71),
    .X(net62),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13225_ (.Y(_06951_),
    .A(\sipo.bit_counter[0] ),
    .B(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13226_ (.B1(_06951_),
    .VDD(VPWR),
    .Y(_00850_),
    .VSS(VGND),
    .A1(\sipo.bit_counter[0] ),
    .A2(_06903_));
 sg13g2_inv_4 _13227_ (.A(net1742),
    .Y(_06952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13228_ (.A(\sipo.word_ready ),
    .B(_06952_),
    .Y(_06953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13229_ (.A(\acc_sum.reg4en.q[0] ),
    .B(_02573_),
    .Y(_06954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13230_ (.A(\acc_sub.reg4en.q[0] ),
    .B(_02576_),
    .Y(_06955_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _13231_ (.A(net1742),
    .B(_02592_),
    .C(_02580_),
    .Y(_06956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _13232_ (.A(_06953_),
    .B(_06954_),
    .C(_06955_),
    .D(_06956_),
    .Y(_06957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13233_ (.B(_02611_),
    .C(_02607_),
    .A(_02600_),
    .Y(_06958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13234_ (.B1(_02592_),
    .VDD(VPWR),
    .Y(_06959_),
    .VSS(VGND),
    .A1(_02598_),
    .A2(_06958_));
 sg13g2_nand2_1 _13235_ (.Y(_06960_),
    .A(net1742),
    .B(\sipo.word_ready ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _13236_ (.Y(_06961_),
    .B(_02628_),
    .A_N(_06960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _13237_ (.X(_06962_),
    .A(_06957_),
    .B(_06959_),
    .C(_06961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13240_ (.Y(_06965_),
    .A(net1711),
    .B(\acc_sub.y[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13241_ (.Y(_06966_),
    .A(net1729),
    .B(\acc_sum.y[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13242_ (.Y(_06967_),
    .A(net1742),
    .B(\sipo.word[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13243_ (.B(_06966_),
    .C(_06967_),
    .A(_06965_),
    .Y(_06968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13244_ (.Y(_06969_),
    .A(net1676),
    .B(_06968_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13245_ (.B1(_06969_),
    .VDD(VPWR),
    .Y(_00849_),
    .VSS(VGND),
    .A1(_01723_),
    .A2(_06962_));
 sg13g2_buf_2 place1728 (.A(_02574_),
    .X(net1728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13247_ (.Y(_06971_),
    .A(_02578_),
    .B(\acc_sub.y[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout92 (.A(net93),
    .X(net92),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13249_ (.Y(_06973_),
    .A(net1729),
    .B(\acc_sum.y[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13250_ (.Y(_06974_),
    .A(net1743),
    .B(\sipo.word[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13251_ (.B(_06973_),
    .C(_06974_),
    .A(_06971_),
    .Y(_06975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _13252_ (.A0(\acc[14] ),
    .A1(_06975_),
    .S(net1676),
    .X(_00848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13254_ (.A(_03244_),
    .B(_02576_),
    .Y(_06977_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13255_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sum.y[13] ),
    .C1(_06977_),
    .B1(net1729),
    .A1(net1743),
    .Y(_06978_),
    .A2(\sipo.word[13] ));
 sg13g2_nor2_1 _13256_ (.A(\acc[13] ),
    .B(net1679),
    .Y(_06979_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13257_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1679),
    .A2(_06978_),
    .Y(_00847_),
    .B1(_06979_));
 sg13g2_inv_2 _13258_ (.Y(_06980_),
    .A(\sipo.word[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _13259_ (.Y(_06981_),
    .B1(\acc_sub.y[12] ),
    .B2(net1711),
    .A2(\acc_sum.y[12] ),
    .A1(net1728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13260_ (.B1(_06981_),
    .VDD(VPWR),
    .Y(_06982_),
    .VSS(VGND),
    .A1(_06980_),
    .A2(_06952_));
 sg13g2_mux2_1 _13261_ (.A0(\acc[12] ),
    .A1(_06982_),
    .S(net1679),
    .X(_00846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13262_ (.A(_03272_),
    .B(_02576_),
    .Y(_06983_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13263_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sum.y[11] ),
    .C1(_06983_),
    .B1(net1729),
    .A1(net1743),
    .Y(_06984_),
    .A2(\sipo.word[11] ));
 sg13g2_nor2_1 _13264_ (.A(\acc[11] ),
    .B(net1679),
    .Y(_06985_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13265_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1679),
    .A2(_06984_),
    .Y(_00845_),
    .B1(_06985_));
 sg13g2_nor2_1 _13266_ (.A(_03283_),
    .B(_02576_),
    .Y(_06986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13267_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sum.y[10] ),
    .C1(_06986_),
    .B1(net1729),
    .A1(net1743),
    .Y(_06987_),
    .A2(\sipo.word[10] ));
 sg13g2_nor2_1 _13268_ (.A(\acc[10] ),
    .B(net1676),
    .Y(_06988_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13269_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1676),
    .A2(_06987_),
    .Y(_00844_),
    .B1(_06988_));
 sg13g2_nor2_1 _13270_ (.A(_03294_),
    .B(_02576_),
    .Y(_06989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13271_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sum.y[9] ),
    .C1(_06989_),
    .B1(net1729),
    .A1(net1743),
    .Y(_06990_),
    .A2(\sipo.word[9] ));
 sg13g2_nor2_1 _13272_ (.A(\acc[9] ),
    .B(net1676),
    .Y(_06991_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13273_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1676),
    .A2(_06990_),
    .Y(_00843_),
    .B1(_06991_));
 sg13g2_nand2_1 _13274_ (.Y(_06992_),
    .A(net1711),
    .B(\acc_sub.y[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13275_ (.Y(_06993_),
    .A(net1729),
    .B(\acc_sum.y[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13276_ (.Y(_06994_),
    .A(net1743),
    .B(\sipo.word[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13277_ (.B(_06993_),
    .C(_06994_),
    .A(_06992_),
    .Y(_06995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _13278_ (.A0(\acc[8] ),
    .A1(_06995_),
    .S(net1678),
    .X(_00842_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13279_ (.A(_03966_),
    .B(_02573_),
    .Y(_06996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13280_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sub.y[7] ),
    .C1(_06996_),
    .B1(_02578_),
    .A1(net1742),
    .Y(_06997_),
    .A2(\sipo.word[7] ));
 sg13g2_nor2_1 _13281_ (.A(\acc[7] ),
    .B(net1676),
    .Y(_06998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13282_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1676),
    .A2(_06997_),
    .Y(_00841_),
    .B1(_06998_));
 sg13g2_inv_2 _13283_ (.Y(_06999_),
    .A(\sipo.word[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13284_ (.A(_06999_),
    .B(_06952_),
    .Y(_07000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13285_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sub.y[6] ),
    .C1(_07000_),
    .B1(_02578_),
    .A1(net1728),
    .Y(_07001_),
    .A2(\acc_sum.y[6] ));
 sg13g2_nor2_1 _13286_ (.A(\acc[6] ),
    .B(net1677),
    .Y(_07002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13287_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1677),
    .A2(_07001_),
    .Y(_00840_),
    .B1(_07002_));
 sg13g2_inv_2 _13288_ (.Y(_07003_),
    .A(\sipo.word[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _13289_ (.Y(_07004_),
    .B1(\acc_sub.y[5] ),
    .B2(net1711),
    .A2(\acc_sum.y[5] ),
    .A1(net1728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13290_ (.B1(_07004_),
    .VDD(VPWR),
    .Y(_07005_),
    .VSS(VGND),
    .A1(_07003_),
    .A2(_06952_));
 sg13g2_mux2_1 _13291_ (.A0(\acc[5] ),
    .A1(_07005_),
    .S(net1679),
    .X(_00839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _13292_ (.Y(_07006_),
    .A(\sipo.word[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13293_ (.A(_07006_),
    .B(_06952_),
    .Y(_07007_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13294_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sub.y[4] ),
    .C1(_07007_),
    .B1(net1711),
    .A1(net1728),
    .Y(_07008_),
    .A2(\acc_sum.y[4] ));
 sg13g2_nor2_1 _13295_ (.A(\acc[4] ),
    .B(net1678),
    .Y(_07009_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13296_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1678),
    .A2(_07008_),
    .Y(_00838_),
    .B1(_07009_));
 sg13g2_inv_2 _13297_ (.Y(_07010_),
    .A(\sipo.word[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13298_ (.A(_07010_),
    .B(_06952_),
    .Y(_07011_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13299_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sub.y[3] ),
    .C1(_07011_),
    .B1(net1711),
    .A1(net1728),
    .Y(_07012_),
    .A2(\acc_sum.y[3] ));
 sg13g2_nor2_1 _13300_ (.A(\acc[3] ),
    .B(net1678),
    .Y(_07013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13301_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1678),
    .A2(_07012_),
    .Y(_00837_),
    .B1(_07013_));
 sg13g2_inv_2 _13302_ (.Y(_07014_),
    .A(\sipo.word[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13303_ (.A(_07014_),
    .B(_06952_),
    .Y(_07015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13304_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sub.y[2] ),
    .C1(_07015_),
    .B1(_02578_),
    .A1(net1728),
    .Y(_07016_),
    .A2(\acc_sum.y[2] ));
 sg13g2_nor2_1 _13305_ (.A(\acc[2] ),
    .B(net1677),
    .Y(_07017_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13306_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1677),
    .A2(_07016_),
    .Y(_00836_),
    .B1(_07017_));
 sg13g2_inv_2 _13307_ (.Y(_07018_),
    .A(\sipo.word[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _13308_ (.A(_07018_),
    .B(_06952_),
    .Y(_07019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _13309_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\acc_sub.y[1] ),
    .C1(_07019_),
    .B1(_02578_),
    .A1(net1728),
    .Y(_07020_),
    .A2(\acc_sum.y[1] ));
 sg13g2_nor2_1 _13310_ (.A(\acc[1] ),
    .B(net1677),
    .Y(_07021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13311_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1677),
    .A2(_07020_),
    .Y(_00835_),
    .B1(_07021_));
 sg13g2_nand2_1 _13312_ (.Y(_07022_),
    .A(_02578_),
    .B(\acc_sub.y[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13313_ (.Y(_07023_),
    .A(net1729),
    .B(\acc_sum.y[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13314_ (.Y(_07024_),
    .A(net1742),
    .B(\sipo.word[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _13315_ (.B(_07023_),
    .C(_07024_),
    .A(_07022_),
    .Y(_07025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _13316_ (.A0(\acc[0] ),
    .A1(_07025_),
    .S(net1678),
    .X(_00834_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _13317_ (.VDD(VPWR),
    .Y(_07026_),
    .A(\sipo.word[15] ),
    .VSS(VGND));
 sg13g2_nand2_2 _13318_ (.Y(_07027_),
    .A(_02563_),
    .B(\sipo.word_ready ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout106 (.A(net107),
    .X(net106),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout105 (.A(net106),
    .X(net105),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout104 (.A(net107),
    .X(net104),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13322_ (.Y(_07031_),
    .A(net1725),
    .B(\fp16_res_pipe.x2[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13323_ (.B1(_07031_),
    .VDD(VPWR),
    .Y(_00833_),
    .VSS(VGND),
    .A1(_07026_),
    .A2(net1725));
 sg13g2_inv_1 _13324_ (.VDD(VPWR),
    .Y(_07032_),
    .A(\sipo.word[14] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13325_ (.Y(_07033_),
    .A(net1725),
    .B(\fp16_res_pipe.x2[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13326_ (.B1(_07033_),
    .VDD(VPWR),
    .Y(_00832_),
    .VSS(VGND),
    .A1(_07032_),
    .A2(net1725));
 sg13g2_inv_1 _13327_ (.VDD(VPWR),
    .Y(_07034_),
    .A(\sipo.word[13] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13328_ (.Y(_07035_),
    .A(net1725),
    .B(\fp16_res_pipe.x2[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13329_ (.B1(_07035_),
    .VDD(VPWR),
    .Y(_00831_),
    .VSS(VGND),
    .A1(_07034_),
    .A2(net1725));
 sg13g2_nand2_1 _13330_ (.Y(_07036_),
    .A(net1724),
    .B(\fp16_res_pipe.x2[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13331_ (.B1(_07036_),
    .VDD(VPWR),
    .Y(_00830_),
    .VSS(VGND),
    .A1(_06980_),
    .A2(net1724));
 sg13g2_inv_1 _13332_ (.VDD(VPWR),
    .Y(_07037_),
    .A(\sipo.word[11] ),
    .VSS(VGND));
 sg13g2_buf_2 fanout103 (.A(net104),
    .X(net103),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13334_ (.Y(_07039_),
    .A(net1726),
    .B(\fp16_res_pipe.x2[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13335_ (.B1(_07039_),
    .VDD(VPWR),
    .Y(_00829_),
    .VSS(VGND),
    .A1(_07037_),
    .A2(net1726));
 sg13g2_inv_1 _13336_ (.VDD(VPWR),
    .Y(_07040_),
    .A(\sipo.word[10] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13337_ (.Y(_07041_),
    .A(net1726),
    .B(\fp16_res_pipe.x2[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13338_ (.B1(_07041_),
    .VDD(VPWR),
    .Y(_00828_),
    .VSS(VGND),
    .A1(_07040_),
    .A2(net1726));
 sg13g2_inv_1 _13339_ (.VDD(VPWR),
    .Y(_07042_),
    .A(\sipo.word[9] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13340_ (.Y(_07043_),
    .A(net1726),
    .B(\fp16_res_pipe.x2[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13341_ (.B1(_07043_),
    .VDD(VPWR),
    .Y(_00827_),
    .VSS(VGND),
    .A1(_07042_),
    .A2(net1726));
 sg13g2_inv_1 _13342_ (.VDD(VPWR),
    .Y(_07044_),
    .A(\sipo.word[8] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13343_ (.Y(_07045_),
    .A(net1726),
    .B(\fp16_res_pipe.x2[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13344_ (.B1(_07045_),
    .VDD(VPWR),
    .Y(_00826_),
    .VSS(VGND),
    .A1(_07044_),
    .A2(net1726));
 sg13g2_inv_1 _13345_ (.VDD(VPWR),
    .Y(_07046_),
    .A(\sipo.word[7] ),
    .VSS(VGND));
 sg13g2_nand2_1 _13346_ (.Y(_07047_),
    .A(_07027_),
    .B(\fp16_res_pipe.x2[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13347_ (.B1(_07047_),
    .VDD(VPWR),
    .Y(_00825_),
    .VSS(VGND),
    .A1(_07046_),
    .A2(_07027_));
 sg13g2_nand2_1 _13348_ (.Y(_07048_),
    .A(net1723),
    .B(\fp16_res_pipe.x2[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13349_ (.B1(_07048_),
    .VDD(VPWR),
    .Y(_00824_),
    .VSS(VGND),
    .A1(_06999_),
    .A2(net1723));
 sg13g2_nand2_1 _13350_ (.Y(_07049_),
    .A(net1724),
    .B(\fp16_res_pipe.x2[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13351_ (.B1(_07049_),
    .VDD(VPWR),
    .Y(_00823_),
    .VSS(VGND),
    .A1(_07003_),
    .A2(net1724));
 sg13g2_nand2_1 _13352_ (.Y(_07050_),
    .A(net1723),
    .B(\fp16_res_pipe.x2[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13353_ (.B1(_07050_),
    .VDD(VPWR),
    .Y(_00822_),
    .VSS(VGND),
    .A1(_07006_),
    .A2(net1723));
 sg13g2_nand2_1 _13354_ (.Y(_07051_),
    .A(net1723),
    .B(\fp16_res_pipe.x2[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13355_ (.B1(_07051_),
    .VDD(VPWR),
    .Y(_00821_),
    .VSS(VGND),
    .A1(_07010_),
    .A2(net1723));
 sg13g2_nand2_1 _13356_ (.Y(_07052_),
    .A(net1724),
    .B(\fp16_res_pipe.x2[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13357_ (.B1(_07052_),
    .VDD(VPWR),
    .Y(_00820_),
    .VSS(VGND),
    .A1(_07014_),
    .A2(net1724));
 sg13g2_nand2_1 _13358_ (.Y(_07053_),
    .A(net1723),
    .B(\fp16_res_pipe.x2[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13359_ (.B1(_07053_),
    .VDD(VPWR),
    .Y(_00819_),
    .VSS(VGND),
    .A1(_07018_),
    .A2(net1723));
 sg13g2_nand2_1 _13360_ (.Y(_07054_),
    .A(_07027_),
    .B(\fp16_res_pipe.x2[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13361_ (.B1(_07054_),
    .VDD(VPWR),
    .Y(_00818_),
    .VSS(VGND),
    .A1(_06941_),
    .A2(_07027_));
 sg13g2_nand2_2 _13362_ (.Y(_07055_),
    .A(_02588_),
    .B(_06960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13366_ (.Y(_07059_),
    .A(net1696),
    .B(\sipo.word[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13367_ (.B1(_07059_),
    .VDD(VPWR),
    .Y(_00817_),
    .VSS(VGND),
    .A1(_03327_),
    .A2(net1696));
 sg13g2_nand2_1 _13368_ (.Y(_07060_),
    .A(net1694),
    .B(\sipo.word[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13369_ (.B1(_07060_),
    .VDD(VPWR),
    .Y(_00816_),
    .VSS(VGND),
    .A1(_05357_),
    .A2(net1694));
 sg13g2_nand2_1 _13370_ (.Y(_07061_),
    .A(net1694),
    .B(\sipo.word[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13371_ (.B1(_07061_),
    .VDD(VPWR),
    .Y(_00815_),
    .VSS(VGND),
    .A1(_05359_),
    .A2(net1694));
 sg13g2_nand2_1 _13372_ (.Y(_07062_),
    .A(net1695),
    .B(\sipo.word[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13373_ (.B1(_07062_),
    .VDD(VPWR),
    .Y(_00814_),
    .VSS(VGND),
    .A1(_06337_),
    .A2(net1694));
 sg13g2_buf_2 fanout141 (.A(net2),
    .X(net141),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13375_ (.Y(_07064_),
    .A(net1695),
    .B(\sipo.word[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13376_ (.B1(_07064_),
    .VDD(VPWR),
    .Y(_00813_),
    .VSS(VGND),
    .A1(_06339_),
    .A2(net1694));
 sg13g2_nand2_1 _13377_ (.Y(_07065_),
    .A(net1695),
    .B(\sipo.word[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13378_ (.B1(_07065_),
    .VDD(VPWR),
    .Y(_00812_),
    .VSS(VGND),
    .A1(_06341_),
    .A2(net1694));
 sg13g2_nand2_1 _13379_ (.Y(_07066_),
    .A(_07055_),
    .B(\sipo.word[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13380_ (.B1(_07066_),
    .VDD(VPWR),
    .Y(_00811_),
    .VSS(VGND),
    .A1(_05367_),
    .A2(_07055_));
 sg13g2_nand2_1 _13381_ (.Y(_07067_),
    .A(net1695),
    .B(\sipo.word[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13382_ (.B1(_07067_),
    .VDD(VPWR),
    .Y(_00810_),
    .VSS(VGND),
    .A1(_03601_),
    .A2(net1695));
 sg13g2_nand2_1 _13383_ (.Y(_07068_),
    .A(net1695),
    .B(\sipo.word[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13384_ (.B1(_07068_),
    .VDD(VPWR),
    .Y(_00809_),
    .VSS(VGND),
    .A1(_03603_),
    .A2(net1695));
 sg13g2_nand2_1 _13385_ (.Y(_07069_),
    .A(net1693),
    .B(\sipo.word[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13386_ (.B1(_07069_),
    .VDD(VPWR),
    .Y(_00808_),
    .VSS(VGND),
    .A1(_06346_),
    .A2(net1694));
 sg13g2_nor2_1 _13387_ (.A(\acc_sub.x2[5] ),
    .B(net1693),
    .Y(_07070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13388_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_07003_),
    .A2(net1695),
    .Y(_00807_),
    .B1(_07070_));
 sg13g2_nor2_1 _13389_ (.A(\acc_sub.x2[4] ),
    .B(net1693),
    .Y(_07071_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13390_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_07006_),
    .A2(net1693),
    .Y(_00806_),
    .B1(_07071_));
 sg13g2_nor2_1 _13391_ (.A(\acc_sub.x2[3] ),
    .B(net1696),
    .Y(_07072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13392_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_07010_),
    .A2(net1696),
    .Y(_00805_),
    .B1(_07072_));
 sg13g2_nor2_1 _13393_ (.A(\acc_sub.x2[2] ),
    .B(net1696),
    .Y(_07073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13394_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_07014_),
    .A2(net1696),
    .Y(_00804_),
    .B1(_07073_));
 sg13g2_nand2_1 _13395_ (.Y(_07074_),
    .A(net1696),
    .B(\sipo.word[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13396_ (.B1(_07074_),
    .VDD(VPWR),
    .Y(_00803_),
    .VSS(VGND),
    .A1(_05382_),
    .A2(net1696));
 sg13g2_nor2_1 _13397_ (.A(\acc_sub.x2[0] ),
    .B(_07055_),
    .Y(_07075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13398_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06941_),
    .A2(_07055_),
    .Y(_00802_),
    .B1(_07075_));
 sg13g2_nand2_2 _13399_ (.Y(_07076_),
    .A(_02566_),
    .B(\sipo.word_ready ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout108 (.A(net113),
    .X(net108),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout107 (.A(net141),
    .X(net107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1916 (.A(net1913),
    .X(net1916),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13403_ (.Y(_07080_),
    .A(net1721),
    .B(\instr[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13404_ (.B1(_07080_),
    .VDD(VPWR),
    .Y(_00801_),
    .VSS(VGND),
    .A1(_07026_),
    .A2(net1721));
 sg13g2_nand2_1 _13405_ (.Y(_07081_),
    .A(net1721),
    .B(\instr[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13406_ (.B1(_07081_),
    .VDD(VPWR),
    .Y(_00800_),
    .VSS(VGND),
    .A1(_07032_),
    .A2(net1721));
 sg13g2_nand2_1 _13407_ (.Y(_07082_),
    .A(net1721),
    .B(\instr[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13408_ (.B1(_07082_),
    .VDD(VPWR),
    .Y(_00799_),
    .VSS(VGND),
    .A1(_07034_),
    .A2(_07076_));
 sg13g2_nand2_1 _13409_ (.Y(_07083_),
    .A(net1721),
    .B(\instr[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13410_ (.B1(_07083_),
    .VDD(VPWR),
    .Y(_00798_),
    .VSS(VGND),
    .A1(_06980_),
    .A2(net1721));
 sg13g2_buf_1 place1918 (.A(net1917),
    .X(net1918),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13412_ (.Y(_07085_),
    .A(net1722),
    .B(\instr[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13413_ (.B1(_07085_),
    .VDD(VPWR),
    .Y(_00797_),
    .VSS(VGND),
    .A1(_07037_),
    .A2(net1722));
 sg13g2_nand2_1 _13414_ (.Y(_07086_),
    .A(net1722),
    .B(\instr[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13415_ (.B1(_07086_),
    .VDD(VPWR),
    .Y(_00796_),
    .VSS(VGND),
    .A1(_07040_),
    .A2(net1722));
 sg13g2_nand2_1 _13416_ (.Y(_07087_),
    .A(net1722),
    .B(\instr[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13417_ (.B1(_07087_),
    .VDD(VPWR),
    .Y(_00795_),
    .VSS(VGND),
    .A1(_07042_),
    .A2(net1722));
 sg13g2_nand2_1 _13418_ (.Y(_07088_),
    .A(net1722),
    .B(\instr[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13419_ (.B1(_07088_),
    .VDD(VPWR),
    .Y(_00794_),
    .VSS(VGND),
    .A1(_07044_),
    .A2(net1722));
 sg13g2_nand2_1 _13420_ (.Y(_07089_),
    .A(net1720),
    .B(\instr[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13421_ (.B1(_07089_),
    .VDD(VPWR),
    .Y(_00793_),
    .VSS(VGND),
    .A1(_07046_),
    .A2(net1720));
 sg13g2_nand2_1 _13422_ (.Y(_07090_),
    .A(net1719),
    .B(\instr[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13423_ (.B1(_07090_),
    .VDD(VPWR),
    .Y(_00792_),
    .VSS(VGND),
    .A1(_06999_),
    .A2(net1719));
 sg13g2_nand2_1 _13424_ (.Y(_07091_),
    .A(net1719),
    .B(\instr[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13425_ (.B1(_07091_),
    .VDD(VPWR),
    .Y(_00791_),
    .VSS(VGND),
    .A1(_07003_),
    .A2(net1719));
 sg13g2_nand2_1 _13426_ (.Y(_07092_),
    .A(net1719),
    .B(\instr[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13427_ (.B1(_07092_),
    .VDD(VPWR),
    .Y(_00790_),
    .VSS(VGND),
    .A1(_07006_),
    .A2(net1719));
 sg13g2_nand2_1 _13428_ (.Y(_07093_),
    .A(net1720),
    .B(\instr[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13429_ (.B1(_07093_),
    .VDD(VPWR),
    .Y(_00789_),
    .VSS(VGND),
    .A1(_07010_),
    .A2(net1719));
 sg13g2_nand2_1 _13430_ (.Y(_07094_),
    .A(_07076_),
    .B(\instr[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13431_ (.B1(_07094_),
    .VDD(VPWR),
    .Y(_00788_),
    .VSS(VGND),
    .A1(_07014_),
    .A2(net1719));
 sg13g2_nand2_1 _13432_ (.Y(_07095_),
    .A(net1720),
    .B(\instr[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13433_ (.B1(_07095_),
    .VDD(VPWR),
    .Y(_00787_),
    .VSS(VGND),
    .A1(_07018_),
    .A2(net1720));
 sg13g2_nand2_1 _13434_ (.Y(_07096_),
    .A(net1720),
    .B(\instr[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13435_ (.B1(_07096_),
    .VDD(VPWR),
    .Y(_00786_),
    .VSS(VGND),
    .A1(_06941_),
    .A2(net1720));
 sg13g2_o21ai_1 _13436_ (.B1(_06906_),
    .VDD(VPWR),
    .Y(_00785_),
    .VSS(VGND),
    .A1(_06911_),
    .A2(_06905_));
 sg13g2_buf_2 fanout61 (.A(net62),
    .X(net61),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13438_ (.Y(_07098_),
    .A(net1752),
    .B(\sipo.shift_reg[14] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13439_ (.B1(_07098_),
    .VDD(VPWR),
    .Y(_00784_),
    .VSS(VGND),
    .A1(_06911_),
    .A2(net1752));
 sg13g2_nand2_1 _13440_ (.Y(_07099_),
    .A(net1751),
    .B(\sipo.shift_reg[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13441_ (.B1(_07099_),
    .VDD(VPWR),
    .Y(_00783_),
    .VSS(VGND),
    .A1(_06914_),
    .A2(net1751));
 sg13g2_nand2_1 _13442_ (.Y(_07100_),
    .A(net1751),
    .B(\sipo.shift_reg[12] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13443_ (.B1(_07100_),
    .VDD(VPWR),
    .Y(_00782_),
    .VSS(VGND),
    .A1(_06916_),
    .A2(net1751));
 sg13g2_nand2_1 _13444_ (.Y(_07101_),
    .A(net1751),
    .B(\sipo.shift_reg[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13445_ (.B1(_07101_),
    .VDD(VPWR),
    .Y(_00781_),
    .VSS(VGND),
    .A1(_06918_),
    .A2(net1751));
 sg13g2_buf_1 fanout60 (.A(net71),
    .X(net60),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _13447_ (.Y(_07103_),
    .A(net1754),
    .B(\sipo.shift_reg[10] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13448_ (.B1(_07103_),
    .VDD(VPWR),
    .Y(_00780_),
    .VSS(VGND),
    .A1(_06920_),
    .A2(net1754));
 sg13g2_nand2_1 _13449_ (.Y(_07104_),
    .A(net1754),
    .B(\sipo.shift_reg[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13450_ (.B1(_07104_),
    .VDD(VPWR),
    .Y(_00779_),
    .VSS(VGND),
    .A1(_06923_),
    .A2(net1754));
 sg13g2_nand2_1 _13451_ (.Y(_07105_),
    .A(net1754),
    .B(\sipo.shift_reg[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13452_ (.B1(_07105_),
    .VDD(VPWR),
    .Y(_00778_),
    .VSS(VGND),
    .A1(_06925_),
    .A2(net1754));
 sg13g2_nand2_1 _13453_ (.Y(_07106_),
    .A(net1754),
    .B(\sipo.shift_reg[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13454_ (.B1(_07106_),
    .VDD(VPWR),
    .Y(_00777_),
    .VSS(VGND),
    .A1(_06927_),
    .A2(net1754));
 sg13g2_nand2_1 _13455_ (.Y(_07107_),
    .A(net1752),
    .B(\sipo.shift_reg[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13456_ (.B1(_07107_),
    .VDD(VPWR),
    .Y(_00776_),
    .VSS(VGND),
    .A1(_06929_),
    .A2(net1752));
 sg13g2_nand2_1 _13457_ (.Y(_07108_),
    .A(net1752),
    .B(\sipo.shift_reg[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13458_ (.B1(_07108_),
    .VDD(VPWR),
    .Y(_00775_),
    .VSS(VGND),
    .A1(_06931_),
    .A2(net1752));
 sg13g2_nand2_1 _13459_ (.Y(_07109_),
    .A(net1752),
    .B(\sipo.shift_reg[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13460_ (.B1(_07109_),
    .VDD(VPWR),
    .Y(_00774_),
    .VSS(VGND),
    .A1(_06933_),
    .A2(net1753));
 sg13g2_nand2_1 _13461_ (.Y(_07110_),
    .A(net1753),
    .B(\sipo.shift_reg[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13462_ (.B1(_07110_),
    .VDD(VPWR),
    .Y(_00773_),
    .VSS(VGND),
    .A1(_06935_),
    .A2(net1753));
 sg13g2_nand2_1 _13463_ (.Y(_07111_),
    .A(net1753),
    .B(\sipo.shift_reg[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13464_ (.B1(_07111_),
    .VDD(VPWR),
    .Y(_00772_),
    .VSS(VGND),
    .A1(_06937_),
    .A2(net1753));
 sg13g2_nand2_1 _13465_ (.Y(_07112_),
    .A(net1753),
    .B(\sipo.shift_reg[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _13466_ (.B1(_07112_),
    .VDD(VPWR),
    .Y(_00771_),
    .VSS(VGND),
    .A1(_06939_),
    .A2(net1753));
 sg13g2_and2_1 _13467_ (.A(_02571_),
    .B(_02564_),
    .X(_00002_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _13468_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06902_),
    .A2(_02582_),
    .Y(_00004_),
    .B1(net1753));
 sg13g2_a21oi_1 _13469_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_06901_),
    .A2(\sipo.receiving ),
    .Y(_00003_),
    .B1(net3));
 sg13g2_inv_1 _13470_ (.VDD(VPWR),
    .Y(_00021_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13471_ (.VDD(VPWR),
    .Y(_00022_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13472_ (.VDD(VPWR),
    .Y(_00023_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13473_ (.VDD(VPWR),
    .Y(_00024_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13474_ (.VDD(VPWR),
    .Y(_00025_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13475_ (.VDD(VPWR),
    .Y(_00026_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13476_ (.VDD(VPWR),
    .Y(_00027_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13477_ (.VDD(VPWR),
    .Y(_00028_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13478_ (.VDD(VPWR),
    .Y(_00029_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13479_ (.VDD(VPWR),
    .Y(_00030_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13480_ (.VDD(VPWR),
    .Y(_00031_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13481_ (.VDD(VPWR),
    .Y(_00032_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13482_ (.VDD(VPWR),
    .Y(_00033_),
    .A(net23),
    .VSS(VGND));
 sg13g2_inv_1 _13483_ (.VDD(VPWR),
    .Y(_00034_),
    .A(net23),
    .VSS(VGND));
 sg13g2_inv_1 _13484_ (.VDD(VPWR),
    .Y(_00035_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _13485_ (.VDD(VPWR),
    .Y(_00036_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13486_ (.VDD(VPWR),
    .Y(_00037_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13487_ (.VDD(VPWR),
    .Y(_00038_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _13488_ (.VDD(VPWR),
    .Y(_00039_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13489_ (.VDD(VPWR),
    .Y(_00040_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _13490_ (.VDD(VPWR),
    .Y(_00041_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13491_ (.VDD(VPWR),
    .Y(_00042_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13492_ (.VDD(VPWR),
    .Y(_00043_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13493_ (.VDD(VPWR),
    .Y(_00044_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13494_ (.VDD(VPWR),
    .Y(_00045_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13495_ (.VDD(VPWR),
    .Y(_00046_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13496_ (.VDD(VPWR),
    .Y(_00047_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13497_ (.VDD(VPWR),
    .Y(_00048_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13498_ (.VDD(VPWR),
    .Y(_00049_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13499_ (.VDD(VPWR),
    .Y(_00050_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13500_ (.VDD(VPWR),
    .Y(_00051_),
    .A(net34),
    .VSS(VGND));
 sg13g2_inv_1 _13501_ (.VDD(VPWR),
    .Y(_00052_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13502_ (.VDD(VPWR),
    .Y(_00053_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _13503_ (.VDD(VPWR),
    .Y(_00054_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _13504_ (.VDD(VPWR),
    .Y(_00055_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13505_ (.VDD(VPWR),
    .Y(_00056_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13506_ (.VDD(VPWR),
    .Y(_00057_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13507_ (.VDD(VPWR),
    .Y(_00058_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13508_ (.VDD(VPWR),
    .Y(_00059_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13509_ (.VDD(VPWR),
    .Y(_00060_),
    .A(net34),
    .VSS(VGND));
 sg13g2_inv_1 _13510_ (.VDD(VPWR),
    .Y(_00061_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13511_ (.VDD(VPWR),
    .Y(_00062_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13512_ (.VDD(VPWR),
    .Y(_00063_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13513_ (.VDD(VPWR),
    .Y(_00064_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13514_ (.VDD(VPWR),
    .Y(_00065_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13515_ (.VDD(VPWR),
    .Y(_00066_),
    .A(net38),
    .VSS(VGND));
 sg13g2_inv_1 _13516_ (.VDD(VPWR),
    .Y(_00067_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _13517_ (.VDD(VPWR),
    .Y(_00068_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13518_ (.VDD(VPWR),
    .Y(_00069_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13519_ (.VDD(VPWR),
    .Y(_00070_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13520_ (.VDD(VPWR),
    .Y(_00071_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13521_ (.VDD(VPWR),
    .Y(_00072_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13522_ (.VDD(VPWR),
    .Y(_00073_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13523_ (.VDD(VPWR),
    .Y(_00074_),
    .A(net86),
    .VSS(VGND));
 sg13g2_inv_1 _13524_ (.VDD(VPWR),
    .Y(_00075_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13525_ (.VDD(VPWR),
    .Y(_00076_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13526_ (.VDD(VPWR),
    .Y(_00077_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13527_ (.VDD(VPWR),
    .Y(_00078_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13528_ (.VDD(VPWR),
    .Y(_00079_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13529_ (.VDD(VPWR),
    .Y(_00080_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13530_ (.VDD(VPWR),
    .Y(_00081_),
    .A(net34),
    .VSS(VGND));
 sg13g2_inv_1 _13531_ (.VDD(VPWR),
    .Y(_00082_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13532_ (.VDD(VPWR),
    .Y(_00083_),
    .A(net37),
    .VSS(VGND));
 sg13g2_inv_1 _13533_ (.VDD(VPWR),
    .Y(_00084_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13534_ (.VDD(VPWR),
    .Y(_00085_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13535_ (.VDD(VPWR),
    .Y(_00086_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13536_ (.VDD(VPWR),
    .Y(_00087_),
    .A(net84),
    .VSS(VGND));
 sg13g2_inv_1 _13537_ (.VDD(VPWR),
    .Y(_00088_),
    .A(net86),
    .VSS(VGND));
 sg13g2_inv_1 _13538_ (.VDD(VPWR),
    .Y(_00089_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _13539_ (.VDD(VPWR),
    .Y(_00090_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _13540_ (.VDD(VPWR),
    .Y(_00091_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _13541_ (.VDD(VPWR),
    .Y(_00092_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _13542_ (.VDD(VPWR),
    .Y(_00093_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _13543_ (.VDD(VPWR),
    .Y(_00094_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13544_ (.VDD(VPWR),
    .Y(_00095_),
    .A(net100),
    .VSS(VGND));
 sg13g2_inv_1 _13545_ (.VDD(VPWR),
    .Y(_00096_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13546_ (.VDD(VPWR),
    .Y(_00097_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _13547_ (.VDD(VPWR),
    .Y(_00098_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13548_ (.VDD(VPWR),
    .Y(_00099_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13549_ (.VDD(VPWR),
    .Y(_00100_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13550_ (.VDD(VPWR),
    .Y(_00101_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13551_ (.VDD(VPWR),
    .Y(_00102_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _13552_ (.VDD(VPWR),
    .Y(_00103_),
    .A(net88),
    .VSS(VGND));
 sg13g2_inv_1 _13553_ (.VDD(VPWR),
    .Y(_00104_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _13554_ (.VDD(VPWR),
    .Y(_00105_),
    .A(net92),
    .VSS(VGND));
 sg13g2_inv_1 _13555_ (.VDD(VPWR),
    .Y(_00106_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _13556_ (.VDD(VPWR),
    .Y(_00107_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13557_ (.VDD(VPWR),
    .Y(_00108_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13558_ (.VDD(VPWR),
    .Y(_00109_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13559_ (.VDD(VPWR),
    .Y(_00110_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13560_ (.VDD(VPWR),
    .Y(_00111_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13561_ (.VDD(VPWR),
    .Y(_00112_),
    .A(net86),
    .VSS(VGND));
 sg13g2_inv_1 _13562_ (.VDD(VPWR),
    .Y(_00113_),
    .A(net83),
    .VSS(VGND));
 sg13g2_inv_1 _13563_ (.VDD(VPWR),
    .Y(_00114_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13564_ (.VDD(VPWR),
    .Y(_00115_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13565_ (.VDD(VPWR),
    .Y(_00116_),
    .A(net82),
    .VSS(VGND));
 sg13g2_inv_1 _13566_ (.VDD(VPWR),
    .Y(_00117_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13567_ (.VDD(VPWR),
    .Y(_00118_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13568_ (.VDD(VPWR),
    .Y(_00119_),
    .A(net33),
    .VSS(VGND));
 sg13g2_inv_1 _13569_ (.VDD(VPWR),
    .Y(_00120_),
    .A(net34),
    .VSS(VGND));
 sg13g2_inv_1 _13570_ (.VDD(VPWR),
    .Y(_00121_),
    .A(net27),
    .VSS(VGND));
 sg13g2_inv_1 _13571_ (.VDD(VPWR),
    .Y(_00122_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13572_ (.VDD(VPWR),
    .Y(_00123_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13573_ (.VDD(VPWR),
    .Y(_00124_),
    .A(net23),
    .VSS(VGND));
 sg13g2_inv_1 _13574_ (.VDD(VPWR),
    .Y(_00125_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13575_ (.VDD(VPWR),
    .Y(_00126_),
    .A(net32),
    .VSS(VGND));
 sg13g2_inv_1 _13576_ (.VDD(VPWR),
    .Y(_00127_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _13577_ (.VDD(VPWR),
    .Y(_00128_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _13578_ (.VDD(VPWR),
    .Y(_00129_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _13579_ (.VDD(VPWR),
    .Y(_00130_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _13580_ (.VDD(VPWR),
    .Y(_00131_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13581_ (.VDD(VPWR),
    .Y(_00132_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _13582_ (.VDD(VPWR),
    .Y(_00133_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13583_ (.VDD(VPWR),
    .Y(_00134_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13584_ (.VDD(VPWR),
    .Y(_00135_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13585_ (.VDD(VPWR),
    .Y(_00136_),
    .A(net115),
    .VSS(VGND));
 sg13g2_inv_1 _13586_ (.VDD(VPWR),
    .Y(_00137_),
    .A(net121),
    .VSS(VGND));
 sg13g2_inv_1 _13587_ (.VDD(VPWR),
    .Y(_00138_),
    .A(net121),
    .VSS(VGND));
 sg13g2_inv_1 _13588_ (.VDD(VPWR),
    .Y(_00139_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _13589_ (.VDD(VPWR),
    .Y(_00140_),
    .A(net121),
    .VSS(VGND));
 sg13g2_inv_1 _13590_ (.VDD(VPWR),
    .Y(_00141_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13591_ (.VDD(VPWR),
    .Y(_00142_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13592_ (.VDD(VPWR),
    .Y(_00143_),
    .A(net121),
    .VSS(VGND));
 sg13g2_inv_1 _13593_ (.VDD(VPWR),
    .Y(_00144_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13594_ (.VDD(VPWR),
    .Y(_00145_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13595_ (.VDD(VPWR),
    .Y(_00146_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13596_ (.VDD(VPWR),
    .Y(_00147_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13597_ (.VDD(VPWR),
    .Y(_00148_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13598_ (.VDD(VPWR),
    .Y(_00149_),
    .A(net62),
    .VSS(VGND));
 sg13g2_inv_1 _13599_ (.VDD(VPWR),
    .Y(_00150_),
    .A(net62),
    .VSS(VGND));
 sg13g2_inv_1 _13600_ (.VDD(VPWR),
    .Y(_00151_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13601_ (.VDD(VPWR),
    .Y(_00152_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13602_ (.VDD(VPWR),
    .Y(_00153_),
    .A(net121),
    .VSS(VGND));
 sg13g2_inv_1 _13603_ (.VDD(VPWR),
    .Y(_00154_),
    .A(net121),
    .VSS(VGND));
 sg13g2_inv_1 _13604_ (.VDD(VPWR),
    .Y(_00155_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13605_ (.VDD(VPWR),
    .Y(_00156_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13606_ (.VDD(VPWR),
    .Y(_00157_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13607_ (.VDD(VPWR),
    .Y(_00158_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13608_ (.VDD(VPWR),
    .Y(_00159_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13609_ (.VDD(VPWR),
    .Y(_00160_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13610_ (.VDD(VPWR),
    .Y(_00161_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13611_ (.VDD(VPWR),
    .Y(_00162_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13612_ (.VDD(VPWR),
    .Y(_00163_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13613_ (.VDD(VPWR),
    .Y(_00164_),
    .A(net112),
    .VSS(VGND));
 sg13g2_inv_1 _13614_ (.VDD(VPWR),
    .Y(_00165_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13615_ (.VDD(VPWR),
    .Y(_00166_),
    .A(net112),
    .VSS(VGND));
 sg13g2_inv_1 _13616_ (.VDD(VPWR),
    .Y(_00167_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13617_ (.VDD(VPWR),
    .Y(_00168_),
    .A(net112),
    .VSS(VGND));
 sg13g2_inv_1 _13618_ (.VDD(VPWR),
    .Y(_00169_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13619_ (.VDD(VPWR),
    .Y(_00170_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13620_ (.VDD(VPWR),
    .Y(_00171_),
    .A(net66),
    .VSS(VGND));
 sg13g2_inv_1 _13621_ (.VDD(VPWR),
    .Y(_00172_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13622_ (.VDD(VPWR),
    .Y(_00173_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13623_ (.VDD(VPWR),
    .Y(_00174_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13624_ (.VDD(VPWR),
    .Y(_00175_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13625_ (.VDD(VPWR),
    .Y(_00176_),
    .A(net69),
    .VSS(VGND));
 sg13g2_inv_1 _13626_ (.VDD(VPWR),
    .Y(_00177_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13627_ (.VDD(VPWR),
    .Y(_00178_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13628_ (.VDD(VPWR),
    .Y(_00179_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13629_ (.VDD(VPWR),
    .Y(_00180_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13630_ (.VDD(VPWR),
    .Y(_00181_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13631_ (.VDD(VPWR),
    .Y(_00182_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13632_ (.VDD(VPWR),
    .Y(_00183_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13633_ (.VDD(VPWR),
    .Y(_00184_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13634_ (.VDD(VPWR),
    .Y(_00185_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13635_ (.VDD(VPWR),
    .Y(_00186_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13636_ (.VDD(VPWR),
    .Y(_00187_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13637_ (.VDD(VPWR),
    .Y(_00188_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _13638_ (.VDD(VPWR),
    .Y(_00189_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _13639_ (.VDD(VPWR),
    .Y(_00190_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _13640_ (.VDD(VPWR),
    .Y(_00191_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13641_ (.VDD(VPWR),
    .Y(_00192_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13642_ (.VDD(VPWR),
    .Y(_00193_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13643_ (.VDD(VPWR),
    .Y(_00194_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13644_ (.VDD(VPWR),
    .Y(_00195_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13645_ (.VDD(VPWR),
    .Y(_00196_),
    .A(net111),
    .VSS(VGND));
 sg13g2_inv_1 _13646_ (.VDD(VPWR),
    .Y(_00197_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13647_ (.VDD(VPWR),
    .Y(_00198_),
    .A(net112),
    .VSS(VGND));
 sg13g2_inv_1 _13648_ (.VDD(VPWR),
    .Y(_00199_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13649_ (.VDD(VPWR),
    .Y(_00200_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13650_ (.VDD(VPWR),
    .Y(_00201_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13651_ (.VDD(VPWR),
    .Y(_00202_),
    .A(net110),
    .VSS(VGND));
 sg13g2_inv_1 _13652_ (.VDD(VPWR),
    .Y(_00203_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13653_ (.VDD(VPWR),
    .Y(_00204_),
    .A(net70),
    .VSS(VGND));
 sg13g2_inv_1 _13654_ (.VDD(VPWR),
    .Y(_00205_),
    .A(net70),
    .VSS(VGND));
 sg13g2_inv_1 _13655_ (.VDD(VPWR),
    .Y(_00206_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13656_ (.VDD(VPWR),
    .Y(_00207_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13657_ (.VDD(VPWR),
    .Y(_00208_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13658_ (.VDD(VPWR),
    .Y(_00209_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13659_ (.VDD(VPWR),
    .Y(_00210_),
    .A(net62),
    .VSS(VGND));
 sg13g2_inv_1 _13660_ (.VDD(VPWR),
    .Y(_00211_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13661_ (.VDD(VPWR),
    .Y(_00212_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13662_ (.VDD(VPWR),
    .Y(_00213_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13663_ (.VDD(VPWR),
    .Y(_00214_),
    .A(net36),
    .VSS(VGND));
 sg13g2_inv_1 _13664_ (.VDD(VPWR),
    .Y(_00215_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13665_ (.VDD(VPWR),
    .Y(_00216_),
    .A(net36),
    .VSS(VGND));
 sg13g2_inv_1 _13666_ (.VDD(VPWR),
    .Y(_00217_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13667_ (.VDD(VPWR),
    .Y(_00218_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13668_ (.VDD(VPWR),
    .Y(_00219_),
    .A(net38),
    .VSS(VGND));
 sg13g2_inv_1 _13669_ (.VDD(VPWR),
    .Y(_00220_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13670_ (.VDD(VPWR),
    .Y(_00221_),
    .A(net122),
    .VSS(VGND));
 sg13g2_inv_1 _13671_ (.VDD(VPWR),
    .Y(_00222_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13672_ (.VDD(VPWR),
    .Y(_00223_),
    .A(net122),
    .VSS(VGND));
 sg13g2_inv_1 _13673_ (.VDD(VPWR),
    .Y(_00224_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13674_ (.VDD(VPWR),
    .Y(_00225_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13675_ (.VDD(VPWR),
    .Y(_00226_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13676_ (.VDD(VPWR),
    .Y(_00227_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13677_ (.VDD(VPWR),
    .Y(_00228_),
    .A(net122),
    .VSS(VGND));
 sg13g2_inv_1 _13678_ (.VDD(VPWR),
    .Y(_00229_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13679_ (.VDD(VPWR),
    .Y(_00230_),
    .A(net120),
    .VSS(VGND));
 sg13g2_inv_1 _13680_ (.VDD(VPWR),
    .Y(_00231_),
    .A(net69),
    .VSS(VGND));
 sg13g2_inv_1 _13681_ (.VDD(VPWR),
    .Y(_00232_),
    .A(net69),
    .VSS(VGND));
 sg13g2_inv_1 _13682_ (.VDD(VPWR),
    .Y(_00233_),
    .A(net69),
    .VSS(VGND));
 sg13g2_inv_1 _13683_ (.VDD(VPWR),
    .Y(_00234_),
    .A(net62),
    .VSS(VGND));
 sg13g2_inv_1 _13684_ (.VDD(VPWR),
    .Y(_00235_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13685_ (.VDD(VPWR),
    .Y(_00236_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13686_ (.VDD(VPWR),
    .Y(_00237_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13687_ (.VDD(VPWR),
    .Y(_00238_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13688_ (.VDD(VPWR),
    .Y(_00239_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13689_ (.VDD(VPWR),
    .Y(_00240_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13690_ (.VDD(VPWR),
    .Y(_00241_),
    .A(net66),
    .VSS(VGND));
 sg13g2_inv_1 _13691_ (.VDD(VPWR),
    .Y(_00242_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13692_ (.VDD(VPWR),
    .Y(_00243_),
    .A(net66),
    .VSS(VGND));
 sg13g2_inv_1 _13693_ (.VDD(VPWR),
    .Y(_00244_),
    .A(net66),
    .VSS(VGND));
 sg13g2_inv_1 _13694_ (.VDD(VPWR),
    .Y(_00245_),
    .A(net66),
    .VSS(VGND));
 sg13g2_inv_1 _13695_ (.VDD(VPWR),
    .Y(_00246_),
    .A(net70),
    .VSS(VGND));
 sg13g2_inv_1 _13696_ (.VDD(VPWR),
    .Y(_00247_),
    .A(net61),
    .VSS(VGND));
 sg13g2_inv_1 _13697_ (.VDD(VPWR),
    .Y(_00248_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13698_ (.VDD(VPWR),
    .Y(_00249_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13699_ (.VDD(VPWR),
    .Y(_00250_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13700_ (.VDD(VPWR),
    .Y(_00251_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13701_ (.VDD(VPWR),
    .Y(_00252_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13702_ (.VDD(VPWR),
    .Y(_00253_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13703_ (.VDD(VPWR),
    .Y(_00254_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13704_ (.VDD(VPWR),
    .Y(_00255_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13705_ (.VDD(VPWR),
    .Y(_00256_),
    .A(net65),
    .VSS(VGND));
 sg13g2_inv_1 _13706_ (.VDD(VPWR),
    .Y(_00257_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13707_ (.VDD(VPWR),
    .Y(_00258_),
    .A(net64),
    .VSS(VGND));
 sg13g2_inv_1 _13708_ (.VDD(VPWR),
    .Y(_00259_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13709_ (.VDD(VPWR),
    .Y(_00260_),
    .A(net64),
    .VSS(VGND));
 sg13g2_inv_1 _13710_ (.VDD(VPWR),
    .Y(_00261_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13711_ (.VDD(VPWR),
    .Y(_00262_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13712_ (.VDD(VPWR),
    .Y(_00263_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _13713_ (.VDD(VPWR),
    .Y(_00264_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _13714_ (.VDD(VPWR),
    .Y(_00265_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _13715_ (.VDD(VPWR),
    .Y(_00266_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13716_ (.VDD(VPWR),
    .Y(_00267_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _13717_ (.VDD(VPWR),
    .Y(_00268_),
    .A(net58),
    .VSS(VGND));
 sg13g2_inv_1 _13718_ (.VDD(VPWR),
    .Y(_00269_),
    .A(net57),
    .VSS(VGND));
 sg13g2_inv_1 _13719_ (.VDD(VPWR),
    .Y(_00270_),
    .A(net60),
    .VSS(VGND));
 sg13g2_inv_1 _13720_ (.VDD(VPWR),
    .Y(_00271_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _13721_ (.VDD(VPWR),
    .Y(_00272_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _13722_ (.VDD(VPWR),
    .Y(_00273_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _13723_ (.VDD(VPWR),
    .Y(_00274_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _13724_ (.VDD(VPWR),
    .Y(_00275_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _13725_ (.VDD(VPWR),
    .Y(_00276_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13726_ (.VDD(VPWR),
    .Y(_00277_),
    .A(net64),
    .VSS(VGND));
 sg13g2_inv_1 _13727_ (.VDD(VPWR),
    .Y(_00278_),
    .A(net64),
    .VSS(VGND));
 sg13g2_inv_1 _13728_ (.VDD(VPWR),
    .Y(_00279_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13729_ (.VDD(VPWR),
    .Y(_00280_),
    .A(net67),
    .VSS(VGND));
 sg13g2_inv_1 _13730_ (.VDD(VPWR),
    .Y(_00281_),
    .A(net64),
    .VSS(VGND));
 sg13g2_inv_1 _13731_ (.VDD(VPWR),
    .Y(_00282_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13732_ (.VDD(VPWR),
    .Y(_00283_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13733_ (.VDD(VPWR),
    .Y(_00284_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13734_ (.VDD(VPWR),
    .Y(_00285_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13735_ (.VDD(VPWR),
    .Y(_00286_),
    .A(net68),
    .VSS(VGND));
 sg13g2_inv_1 _13736_ (.VDD(VPWR),
    .Y(_00287_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13737_ (.VDD(VPWR),
    .Y(_00288_),
    .A(net55),
    .VSS(VGND));
 sg13g2_inv_1 _13738_ (.VDD(VPWR),
    .Y(_00289_),
    .A(net63),
    .VSS(VGND));
 sg13g2_inv_1 _13739_ (.VDD(VPWR),
    .Y(_00290_),
    .A(net55),
    .VSS(VGND));
 sg13g2_inv_1 _13740_ (.VDD(VPWR),
    .Y(_00291_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _13741_ (.VDD(VPWR),
    .Y(_00292_),
    .A(net86),
    .VSS(VGND));
 sg13g2_inv_1 _13742_ (.VDD(VPWR),
    .Y(_00293_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _13743_ (.VDD(VPWR),
    .Y(_00294_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13744_ (.VDD(VPWR),
    .Y(_00295_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _13745_ (.VDD(VPWR),
    .Y(_00296_),
    .A(net118),
    .VSS(VGND));
 sg13g2_inv_1 _13746_ (.VDD(VPWR),
    .Y(_00297_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13747_ (.VDD(VPWR),
    .Y(_00298_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _13748_ (.VDD(VPWR),
    .Y(_00299_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13749_ (.VDD(VPWR),
    .Y(_00300_),
    .A(net123),
    .VSS(VGND));
 sg13g2_inv_1 _13750_ (.VDD(VPWR),
    .Y(_00301_),
    .A(net115),
    .VSS(VGND));
 sg13g2_inv_1 _13751_ (.VDD(VPWR),
    .Y(_00302_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _13752_ (.VDD(VPWR),
    .Y(_00303_),
    .A(net109),
    .VSS(VGND));
 sg13g2_inv_1 _13753_ (.VDD(VPWR),
    .Y(_00304_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13754_ (.VDD(VPWR),
    .Y(_00305_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13755_ (.VDD(VPWR),
    .Y(_00306_),
    .A(net85),
    .VSS(VGND));
 sg13g2_inv_1 _13756_ (.VDD(VPWR),
    .Y(_00307_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13757_ (.VDD(VPWR),
    .Y(_00308_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13758_ (.VDD(VPWR),
    .Y(_00309_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13759_ (.VDD(VPWR),
    .Y(_00310_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _13760_ (.VDD(VPWR),
    .Y(_00311_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _13761_ (.VDD(VPWR),
    .Y(_00312_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _13762_ (.VDD(VPWR),
    .Y(_00313_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _13763_ (.VDD(VPWR),
    .Y(_00314_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _13764_ (.VDD(VPWR),
    .Y(_00315_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _13765_ (.VDD(VPWR),
    .Y(_00316_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _13766_ (.VDD(VPWR),
    .Y(_00317_),
    .A(net115),
    .VSS(VGND));
 sg13g2_inv_1 _13767_ (.VDD(VPWR),
    .Y(_00318_),
    .A(net59),
    .VSS(VGND));
 sg13g2_inv_1 _13768_ (.VDD(VPWR),
    .Y(_00319_),
    .A(net109),
    .VSS(VGND));
 sg13g2_inv_1 _13769_ (.VDD(VPWR),
    .Y(_00320_),
    .A(net109),
    .VSS(VGND));
 sg13g2_inv_1 _13770_ (.VDD(VPWR),
    .Y(_00321_),
    .A(net109),
    .VSS(VGND));
 sg13g2_inv_1 _13771_ (.VDD(VPWR),
    .Y(_00322_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13772_ (.VDD(VPWR),
    .Y(_00323_),
    .A(net38),
    .VSS(VGND));
 sg13g2_inv_1 _13773_ (.VDD(VPWR),
    .Y(_00324_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13774_ (.VDD(VPWR),
    .Y(_00325_),
    .A(net108),
    .VSS(VGND));
 sg13g2_inv_1 _13775_ (.VDD(VPWR),
    .Y(_00326_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _13776_ (.VDD(VPWR),
    .Y(_00327_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _13777_ (.VDD(VPWR),
    .Y(_00328_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _13778_ (.VDD(VPWR),
    .Y(_00329_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13779_ (.VDD(VPWR),
    .Y(_00330_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _13780_ (.VDD(VPWR),
    .Y(_00331_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _13781_ (.VDD(VPWR),
    .Y(_00332_),
    .A(net126),
    .VSS(VGND));
 sg13g2_inv_1 _13782_ (.VDD(VPWR),
    .Y(_00333_),
    .A(net126),
    .VSS(VGND));
 sg13g2_inv_1 _13783_ (.VDD(VPWR),
    .Y(_00334_),
    .A(net125),
    .VSS(VGND));
 sg13g2_inv_1 _13784_ (.VDD(VPWR),
    .Y(_00335_),
    .A(net126),
    .VSS(VGND));
 sg13g2_inv_1 _13785_ (.VDD(VPWR),
    .Y(_00336_),
    .A(net126),
    .VSS(VGND));
 sg13g2_inv_1 _13786_ (.VDD(VPWR),
    .Y(_00337_),
    .A(net126),
    .VSS(VGND));
 sg13g2_inv_1 _13787_ (.VDD(VPWR),
    .Y(_00338_),
    .A(net74),
    .VSS(VGND));
 sg13g2_inv_1 _13788_ (.VDD(VPWR),
    .Y(_00339_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _13789_ (.VDD(VPWR),
    .Y(_00340_),
    .A(net74),
    .VSS(VGND));
 sg13g2_inv_1 _13790_ (.VDD(VPWR),
    .Y(_00341_),
    .A(net20),
    .VSS(VGND));
 sg13g2_inv_1 _13791_ (.VDD(VPWR),
    .Y(_00342_),
    .A(net20),
    .VSS(VGND));
 sg13g2_inv_1 _13792_ (.VDD(VPWR),
    .Y(_00343_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _13793_ (.VDD(VPWR),
    .Y(_00344_),
    .A(net74),
    .VSS(VGND));
 sg13g2_inv_1 _13794_ (.VDD(VPWR),
    .Y(_00345_),
    .A(net20),
    .VSS(VGND));
 sg13g2_inv_1 _13795_ (.VDD(VPWR),
    .Y(_00346_),
    .A(net20),
    .VSS(VGND));
 sg13g2_inv_1 _13796_ (.VDD(VPWR),
    .Y(_00347_),
    .A(net20),
    .VSS(VGND));
 sg13g2_inv_1 _13797_ (.VDD(VPWR),
    .Y(_00348_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _13798_ (.VDD(VPWR),
    .Y(_00349_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13799_ (.VDD(VPWR),
    .Y(_00350_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13800_ (.VDD(VPWR),
    .Y(_00351_),
    .A(net74),
    .VSS(VGND));
 sg13g2_inv_1 _13801_ (.VDD(VPWR),
    .Y(_00352_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13802_ (.VDD(VPWR),
    .Y(_00353_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13803_ (.VDD(VPWR),
    .Y(_00354_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _13804_ (.VDD(VPWR),
    .Y(_00355_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13805_ (.VDD(VPWR),
    .Y(_00356_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13806_ (.VDD(VPWR),
    .Y(_00357_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _13807_ (.VDD(VPWR),
    .Y(_00358_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _13808_ (.VDD(VPWR),
    .Y(_00359_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _13809_ (.VDD(VPWR),
    .Y(_00360_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _13810_ (.VDD(VPWR),
    .Y(_00361_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _13811_ (.VDD(VPWR),
    .Y(_00362_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _13812_ (.VDD(VPWR),
    .Y(_00363_),
    .A(net78),
    .VSS(VGND));
 sg13g2_inv_1 _13813_ (.VDD(VPWR),
    .Y(_00364_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _13814_ (.VDD(VPWR),
    .Y(_00365_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _13815_ (.VDD(VPWR),
    .Y(_00366_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _13816_ (.VDD(VPWR),
    .Y(_00367_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _13817_ (.VDD(VPWR),
    .Y(_00368_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _13818_ (.VDD(VPWR),
    .Y(_00369_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _13819_ (.VDD(VPWR),
    .Y(_00370_),
    .A(net62),
    .VSS(VGND));
 sg13g2_inv_1 _13820_ (.VDD(VPWR),
    .Y(_00371_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _13821_ (.VDD(VPWR),
    .Y(_00372_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _13822_ (.VDD(VPWR),
    .Y(_00373_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _13823_ (.VDD(VPWR),
    .Y(_00374_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _13824_ (.VDD(VPWR),
    .Y(_00375_),
    .A(net14),
    .VSS(VGND));
 sg13g2_inv_1 _13825_ (.VDD(VPWR),
    .Y(_00376_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13826_ (.VDD(VPWR),
    .Y(_00377_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13827_ (.VDD(VPWR),
    .Y(_00378_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13828_ (.VDD(VPWR),
    .Y(_00379_),
    .A(net47),
    .VSS(VGND));
 sg13g2_inv_1 _13829_ (.VDD(VPWR),
    .Y(_00380_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13830_ (.VDD(VPWR),
    .Y(_00381_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13831_ (.VDD(VPWR),
    .Y(_00382_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13832_ (.VDD(VPWR),
    .Y(_00383_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _13833_ (.VDD(VPWR),
    .Y(_00384_),
    .A(net56),
    .VSS(VGND));
 sg13g2_inv_1 _13834_ (.VDD(VPWR),
    .Y(_00385_),
    .A(net14),
    .VSS(VGND));
 sg13g2_inv_1 _13835_ (.VDD(VPWR),
    .Y(_00386_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13836_ (.VDD(VPWR),
    .Y(_00387_),
    .A(net14),
    .VSS(VGND));
 sg13g2_inv_1 _13837_ (.VDD(VPWR),
    .Y(_00388_),
    .A(net14),
    .VSS(VGND));
 sg13g2_inv_1 _13838_ (.VDD(VPWR),
    .Y(_00389_),
    .A(net54),
    .VSS(VGND));
 sg13g2_inv_1 _13839_ (.VDD(VPWR),
    .Y(_00390_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13840_ (.VDD(VPWR),
    .Y(_00391_),
    .A(net36),
    .VSS(VGND));
 sg13g2_inv_1 _13841_ (.VDD(VPWR),
    .Y(_00392_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13842_ (.VDD(VPWR),
    .Y(_00393_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13843_ (.VDD(VPWR),
    .Y(_00394_),
    .A(net36),
    .VSS(VGND));
 sg13g2_inv_1 _13844_ (.VDD(VPWR),
    .Y(_00395_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _13845_ (.VDD(VPWR),
    .Y(_00396_),
    .A(net31),
    .VSS(VGND));
 sg13g2_inv_1 _13846_ (.VDD(VPWR),
    .Y(_00397_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13847_ (.VDD(VPWR),
    .Y(_00398_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13848_ (.VDD(VPWR),
    .Y(_00399_),
    .A(net31),
    .VSS(VGND));
 sg13g2_inv_1 _13849_ (.VDD(VPWR),
    .Y(_00400_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _13850_ (.VDD(VPWR),
    .Y(_00401_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13851_ (.VDD(VPWR),
    .Y(_00402_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _13852_ (.VDD(VPWR),
    .Y(_00403_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _13853_ (.VDD(VPWR),
    .Y(_00404_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _13854_ (.VDD(VPWR),
    .Y(_00405_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13855_ (.VDD(VPWR),
    .Y(_00406_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _13856_ (.VDD(VPWR),
    .Y(_00407_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _13857_ (.VDD(VPWR),
    .Y(_00408_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _13858_ (.VDD(VPWR),
    .Y(_00409_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _13859_ (.VDD(VPWR),
    .Y(_00410_),
    .A(net14),
    .VSS(VGND));
 sg13g2_inv_1 _13860_ (.VDD(VPWR),
    .Y(_00411_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _13861_ (.VDD(VPWR),
    .Y(_00412_),
    .A(net47),
    .VSS(VGND));
 sg13g2_inv_1 _13862_ (.VDD(VPWR),
    .Y(_00413_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13863_ (.VDD(VPWR),
    .Y(_00414_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13864_ (.VDD(VPWR),
    .Y(_00415_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _13865_ (.VDD(VPWR),
    .Y(_00416_),
    .A(net56),
    .VSS(VGND));
 sg13g2_inv_1 _13866_ (.VDD(VPWR),
    .Y(_00417_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13867_ (.VDD(VPWR),
    .Y(_00418_),
    .A(net51),
    .VSS(VGND));
 sg13g2_inv_1 _13868_ (.VDD(VPWR),
    .Y(_00419_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13869_ (.VDD(VPWR),
    .Y(_00420_),
    .A(net14),
    .VSS(VGND));
 sg13g2_inv_1 _13870_ (.VDD(VPWR),
    .Y(_00421_),
    .A(net50),
    .VSS(VGND));
 sg13g2_inv_1 _13871_ (.VDD(VPWR),
    .Y(_00422_),
    .A(net45),
    .VSS(VGND));
 sg13g2_inv_1 _13872_ (.VDD(VPWR),
    .Y(_00423_),
    .A(net45),
    .VSS(VGND));
 sg13g2_inv_1 _13873_ (.VDD(VPWR),
    .Y(_00424_),
    .A(net45),
    .VSS(VGND));
 sg13g2_inv_1 _13874_ (.VDD(VPWR),
    .Y(_00425_),
    .A(net45),
    .VSS(VGND));
 sg13g2_inv_1 _13875_ (.VDD(VPWR),
    .Y(_00426_),
    .A(net53),
    .VSS(VGND));
 sg13g2_inv_1 _13876_ (.VDD(VPWR),
    .Y(_00427_),
    .A(net53),
    .VSS(VGND));
 sg13g2_inv_1 _13877_ (.VDD(VPWR),
    .Y(_00428_),
    .A(net53),
    .VSS(VGND));
 sg13g2_inv_1 _13878_ (.VDD(VPWR),
    .Y(_00429_),
    .A(net53),
    .VSS(VGND));
 sg13g2_inv_1 _13879_ (.VDD(VPWR),
    .Y(_00430_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13880_ (.VDD(VPWR),
    .Y(_00431_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13881_ (.VDD(VPWR),
    .Y(_00432_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13882_ (.VDD(VPWR),
    .Y(_00433_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13883_ (.VDD(VPWR),
    .Y(_00434_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13884_ (.VDD(VPWR),
    .Y(_00435_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13885_ (.VDD(VPWR),
    .Y(_00436_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13886_ (.VDD(VPWR),
    .Y(_00437_),
    .A(net48),
    .VSS(VGND));
 sg13g2_inv_1 _13887_ (.VDD(VPWR),
    .Y(_00438_),
    .A(net49),
    .VSS(VGND));
 sg13g2_inv_1 _13888_ (.VDD(VPWR),
    .Y(_00439_),
    .A(net49),
    .VSS(VGND));
 sg13g2_inv_1 _13889_ (.VDD(VPWR),
    .Y(_00440_),
    .A(net49),
    .VSS(VGND));
 sg13g2_inv_1 _13890_ (.VDD(VPWR),
    .Y(_00441_),
    .A(net49),
    .VSS(VGND));
 sg13g2_inv_1 _13891_ (.VDD(VPWR),
    .Y(_00442_),
    .A(net53),
    .VSS(VGND));
 sg13g2_inv_1 _13892_ (.VDD(VPWR),
    .Y(_00443_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _13893_ (.VDD(VPWR),
    .Y(_00444_),
    .A(net35),
    .VSS(VGND));
 sg13g2_inv_1 _13894_ (.VDD(VPWR),
    .Y(_00445_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _13895_ (.VDD(VPWR),
    .Y(_00446_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13896_ (.VDD(VPWR),
    .Y(_00447_),
    .A(net17),
    .VSS(VGND));
 sg13g2_inv_1 _13897_ (.VDD(VPWR),
    .Y(_00448_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13898_ (.VDD(VPWR),
    .Y(_00449_),
    .A(net17),
    .VSS(VGND));
 sg13g2_inv_1 _13899_ (.VDD(VPWR),
    .Y(_00450_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13900_ (.VDD(VPWR),
    .Y(_00451_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13901_ (.VDD(VPWR),
    .Y(_00452_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13902_ (.VDD(VPWR),
    .Y(_00453_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13903_ (.VDD(VPWR),
    .Y(_00454_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13904_ (.VDD(VPWR),
    .Y(_00455_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13905_ (.VDD(VPWR),
    .Y(_00456_),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _13906_ (.VDD(VPWR),
    .Y(_00457_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13907_ (.VDD(VPWR),
    .Y(_00458_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13908_ (.VDD(VPWR),
    .Y(_00459_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13909_ (.VDD(VPWR),
    .Y(_00460_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13910_ (.VDD(VPWR),
    .Y(_00461_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13911_ (.VDD(VPWR),
    .Y(_00462_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13912_ (.VDD(VPWR),
    .Y(_00463_),
    .A(net27),
    .VSS(VGND));
 sg13g2_inv_1 _13913_ (.VDD(VPWR),
    .Y(_00464_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13914_ (.VDD(VPWR),
    .Y(_00465_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13915_ (.VDD(VPWR),
    .Y(_00466_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13916_ (.VDD(VPWR),
    .Y(_00467_),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _13917_ (.VDD(VPWR),
    .Y(_00468_),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _13918_ (.VDD(VPWR),
    .Y(_00469_),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _13919_ (.VDD(VPWR),
    .Y(_00470_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13920_ (.VDD(VPWR),
    .Y(_00471_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13921_ (.VDD(VPWR),
    .Y(_00472_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13922_ (.VDD(VPWR),
    .Y(_00473_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13923_ (.VDD(VPWR),
    .Y(_00474_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13924_ (.VDD(VPWR),
    .Y(_00475_),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 _13925_ (.VDD(VPWR),
    .Y(_00476_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13926_ (.VDD(VPWR),
    .Y(_00477_),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 _13927_ (.VDD(VPWR),
    .Y(_00478_),
    .A(net8),
    .VSS(VGND));
 sg13g2_inv_1 _13928_ (.VDD(VPWR),
    .Y(_00479_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13929_ (.VDD(VPWR),
    .Y(_00480_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13930_ (.VDD(VPWR),
    .Y(_00481_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13931_ (.VDD(VPWR),
    .Y(_00482_),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 _13932_ (.VDD(VPWR),
    .Y(_00483_),
    .A(net5),
    .VSS(VGND));
 sg13g2_inv_1 _13933_ (.VDD(VPWR),
    .Y(_00484_),
    .A(net6),
    .VSS(VGND));
 sg13g2_inv_1 _13934_ (.VDD(VPWR),
    .Y(_00485_),
    .A(net11),
    .VSS(VGND));
 sg13g2_inv_1 _13935_ (.VDD(VPWR),
    .Y(_00486_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13936_ (.VDD(VPWR),
    .Y(_00487_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13937_ (.VDD(VPWR),
    .Y(_00488_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13938_ (.VDD(VPWR),
    .Y(_00489_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13939_ (.VDD(VPWR),
    .Y(_00490_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13940_ (.VDD(VPWR),
    .Y(_00491_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13941_ (.VDD(VPWR),
    .Y(_00492_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13942_ (.VDD(VPWR),
    .Y(_00493_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13943_ (.VDD(VPWR),
    .Y(_00494_),
    .A(net27),
    .VSS(VGND));
 sg13g2_inv_1 _13944_ (.VDD(VPWR),
    .Y(_00495_),
    .A(net27),
    .VSS(VGND));
 sg13g2_inv_1 _13945_ (.VDD(VPWR),
    .Y(_00496_),
    .A(net27),
    .VSS(VGND));
 sg13g2_inv_1 _13946_ (.VDD(VPWR),
    .Y(_00497_),
    .A(net29),
    .VSS(VGND));
 sg13g2_inv_1 _13947_ (.VDD(VPWR),
    .Y(_00498_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13948_ (.VDD(VPWR),
    .Y(_00499_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13949_ (.VDD(VPWR),
    .Y(_00500_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13950_ (.VDD(VPWR),
    .Y(_00501_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13951_ (.VDD(VPWR),
    .Y(_00502_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _13952_ (.VDD(VPWR),
    .Y(_00503_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _13953_ (.VDD(VPWR),
    .Y(_00504_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13954_ (.VDD(VPWR),
    .Y(_00505_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _13955_ (.VDD(VPWR),
    .Y(_00506_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13956_ (.VDD(VPWR),
    .Y(_00507_),
    .A(net92),
    .VSS(VGND));
 sg13g2_inv_1 _13957_ (.VDD(VPWR),
    .Y(_00508_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _13958_ (.VDD(VPWR),
    .Y(_00509_),
    .A(net96),
    .VSS(VGND));
 sg13g2_inv_1 _13959_ (.VDD(VPWR),
    .Y(_00510_),
    .A(net96),
    .VSS(VGND));
 sg13g2_inv_1 _13960_ (.VDD(VPWR),
    .Y(_00511_),
    .A(net96),
    .VSS(VGND));
 sg13g2_inv_1 _13961_ (.VDD(VPWR),
    .Y(_00512_),
    .A(net97),
    .VSS(VGND));
 sg13g2_inv_1 _13962_ (.VDD(VPWR),
    .Y(_00513_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _13963_ (.VDD(VPWR),
    .Y(_00514_),
    .A(net18),
    .VSS(VGND));
 sg13g2_inv_1 _13964_ (.VDD(VPWR),
    .Y(_00515_),
    .A(net18),
    .VSS(VGND));
 sg13g2_inv_1 _13965_ (.VDD(VPWR),
    .Y(_00516_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13966_ (.VDD(VPWR),
    .Y(_00517_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13967_ (.VDD(VPWR),
    .Y(_00518_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13968_ (.VDD(VPWR),
    .Y(_00519_),
    .A(net7),
    .VSS(VGND));
 sg13g2_inv_1 _13969_ (.VDD(VPWR),
    .Y(_00520_),
    .A(net18),
    .VSS(VGND));
 sg13g2_inv_1 _13970_ (.VDD(VPWR),
    .Y(_00521_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13971_ (.VDD(VPWR),
    .Y(_00522_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13972_ (.VDD(VPWR),
    .Y(_00523_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13973_ (.VDD(VPWR),
    .Y(_00524_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13974_ (.VDD(VPWR),
    .Y(_00525_),
    .A(net17),
    .VSS(VGND));
 sg13g2_inv_1 _13975_ (.VDD(VPWR),
    .Y(_00526_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13976_ (.VDD(VPWR),
    .Y(_00527_),
    .A(net17),
    .VSS(VGND));
 sg13g2_inv_1 _13977_ (.VDD(VPWR),
    .Y(_00528_),
    .A(net16),
    .VSS(VGND));
 sg13g2_inv_1 _13978_ (.VDD(VPWR),
    .Y(_00529_),
    .A(net26),
    .VSS(VGND));
 sg13g2_inv_1 _13979_ (.VDD(VPWR),
    .Y(_00530_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13980_ (.VDD(VPWR),
    .Y(_00531_),
    .A(net13),
    .VSS(VGND));
 sg13g2_inv_1 _13981_ (.VDD(VPWR),
    .Y(_00532_),
    .A(net12),
    .VSS(VGND));
 sg13g2_inv_1 _13982_ (.VDD(VPWR),
    .Y(_00533_),
    .A(net13),
    .VSS(VGND));
 sg13g2_inv_1 _13983_ (.VDD(VPWR),
    .Y(_00534_),
    .A(net13),
    .VSS(VGND));
 sg13g2_inv_1 _13984_ (.VDD(VPWR),
    .Y(_00535_),
    .A(net25),
    .VSS(VGND));
 sg13g2_inv_1 _13985_ (.VDD(VPWR),
    .Y(_00536_),
    .A(net28),
    .VSS(VGND));
 sg13g2_inv_1 _13986_ (.VDD(VPWR),
    .Y(_00537_),
    .A(net28),
    .VSS(VGND));
 sg13g2_inv_1 _13987_ (.VDD(VPWR),
    .Y(_00538_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13988_ (.VDD(VPWR),
    .Y(_00539_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13989_ (.VDD(VPWR),
    .Y(_00540_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13990_ (.VDD(VPWR),
    .Y(_00541_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13991_ (.VDD(VPWR),
    .Y(_00542_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13992_ (.VDD(VPWR),
    .Y(_00543_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13993_ (.VDD(VPWR),
    .Y(_00544_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13994_ (.VDD(VPWR),
    .Y(_00545_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13995_ (.VDD(VPWR),
    .Y(_00546_),
    .A(net15),
    .VSS(VGND));
 sg13g2_inv_1 _13996_ (.VDD(VPWR),
    .Y(_00547_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13997_ (.VDD(VPWR),
    .Y(_00548_),
    .A(net10),
    .VSS(VGND));
 sg13g2_inv_1 _13998_ (.VDD(VPWR),
    .Y(_00549_),
    .A(net9),
    .VSS(VGND));
 sg13g2_inv_1 _13999_ (.VDD(VPWR),
    .Y(_00550_),
    .A(net30),
    .VSS(VGND));
 sg13g2_inv_1 _14000_ (.VDD(VPWR),
    .Y(_00551_),
    .A(net13),
    .VSS(VGND));
 sg13g2_inv_1 _14001_ (.VDD(VPWR),
    .Y(_00552_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _14002_ (.VDD(VPWR),
    .Y(_00553_),
    .A(net78),
    .VSS(VGND));
 sg13g2_inv_1 _14003_ (.VDD(VPWR),
    .Y(_00554_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _14004_ (.VDD(VPWR),
    .Y(_00555_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _14005_ (.VDD(VPWR),
    .Y(_00556_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _14006_ (.VDD(VPWR),
    .Y(_00557_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _14007_ (.VDD(VPWR),
    .Y(_00558_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _14008_ (.VDD(VPWR),
    .Y(_00559_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _14009_ (.VDD(VPWR),
    .Y(_00560_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _14010_ (.VDD(VPWR),
    .Y(_00561_),
    .A(net19),
    .VSS(VGND));
 sg13g2_inv_1 _14011_ (.VDD(VPWR),
    .Y(_00562_),
    .A(net21),
    .VSS(VGND));
 sg13g2_inv_1 _14012_ (.VDD(VPWR),
    .Y(_00563_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _14013_ (.VDD(VPWR),
    .Y(_00564_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _14014_ (.VDD(VPWR),
    .Y(_00565_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _14015_ (.VDD(VPWR),
    .Y(_00566_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _14016_ (.VDD(VPWR),
    .Y(_00567_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _14017_ (.VDD(VPWR),
    .Y(_00568_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _14018_ (.VDD(VPWR),
    .Y(_00569_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _14019_ (.VDD(VPWR),
    .Y(_00570_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _14020_ (.VDD(VPWR),
    .Y(_00571_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _14021_ (.VDD(VPWR),
    .Y(_00572_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _14022_ (.VDD(VPWR),
    .Y(_00573_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _14023_ (.VDD(VPWR),
    .Y(_00574_),
    .A(net100),
    .VSS(VGND));
 sg13g2_inv_1 _14024_ (.VDD(VPWR),
    .Y(_00575_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _14025_ (.VDD(VPWR),
    .Y(_00576_),
    .A(net100),
    .VSS(VGND));
 sg13g2_inv_1 _14026_ (.VDD(VPWR),
    .Y(_00577_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _14027_ (.VDD(VPWR),
    .Y(_00578_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14028_ (.VDD(VPWR),
    .Y(_00579_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _14029_ (.VDD(VPWR),
    .Y(_00580_),
    .A(net99),
    .VSS(VGND));
 sg13g2_inv_1 _14030_ (.VDD(VPWR),
    .Y(_00581_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _14031_ (.VDD(VPWR),
    .Y(_00582_),
    .A(net106),
    .VSS(VGND));
 sg13g2_inv_1 _14032_ (.VDD(VPWR),
    .Y(_00583_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _14033_ (.VDD(VPWR),
    .Y(_00584_),
    .A(net98),
    .VSS(VGND));
 sg13g2_inv_1 _14034_ (.VDD(VPWR),
    .Y(_00585_),
    .A(net107),
    .VSS(VGND));
 sg13g2_inv_1 _14035_ (.VDD(VPWR),
    .Y(_00586_),
    .A(net106),
    .VSS(VGND));
 sg13g2_inv_1 _14036_ (.VDD(VPWR),
    .Y(_00587_),
    .A(net99),
    .VSS(VGND));
 sg13g2_inv_1 _14037_ (.VDD(VPWR),
    .Y(_00588_),
    .A(net73),
    .VSS(VGND));
 sg13g2_inv_1 _14038_ (.VDD(VPWR),
    .Y(_00589_),
    .A(net77),
    .VSS(VGND));
 sg13g2_inv_1 _14039_ (.VDD(VPWR),
    .Y(_00590_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _14040_ (.VDD(VPWR),
    .Y(_00591_),
    .A(net74),
    .VSS(VGND));
 sg13g2_inv_1 _14041_ (.VDD(VPWR),
    .Y(_00592_),
    .A(net76),
    .VSS(VGND));
 sg13g2_inv_1 _14042_ (.VDD(VPWR),
    .Y(_00593_),
    .A(net20),
    .VSS(VGND));
 sg13g2_inv_1 _14043_ (.VDD(VPWR),
    .Y(_00594_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _14044_ (.VDD(VPWR),
    .Y(_00595_),
    .A(net78),
    .VSS(VGND));
 sg13g2_inv_1 _14045_ (.VDD(VPWR),
    .Y(_00596_),
    .A(net76),
    .VSS(VGND));
 sg13g2_inv_1 _14046_ (.VDD(VPWR),
    .Y(_00597_),
    .A(net86),
    .VSS(VGND));
 sg13g2_inv_1 _14047_ (.VDD(VPWR),
    .Y(_00598_),
    .A(net76),
    .VSS(VGND));
 sg13g2_inv_1 _14048_ (.VDD(VPWR),
    .Y(_00599_),
    .A(net75),
    .VSS(VGND));
 sg13g2_inv_1 _14049_ (.VDD(VPWR),
    .Y(_00600_),
    .A(net23),
    .VSS(VGND));
 sg13g2_inv_1 _14050_ (.VDD(VPWR),
    .Y(_00601_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _14051_ (.VDD(VPWR),
    .Y(_00602_),
    .A(net22),
    .VSS(VGND));
 sg13g2_inv_1 _14052_ (.VDD(VPWR),
    .Y(_00603_),
    .A(net87),
    .VSS(VGND));
 sg13g2_inv_1 _14053_ (.VDD(VPWR),
    .Y(_00604_),
    .A(net81),
    .VSS(VGND));
 sg13g2_inv_1 _14054_ (.VDD(VPWR),
    .Y(_00605_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _14055_ (.VDD(VPWR),
    .Y(_00606_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _14056_ (.VDD(VPWR),
    .Y(_00607_),
    .A(net96),
    .VSS(VGND));
 sg13g2_inv_1 _14057_ (.VDD(VPWR),
    .Y(_00608_),
    .A(net78),
    .VSS(VGND));
 sg13g2_inv_1 _14058_ (.VDD(VPWR),
    .Y(_00609_),
    .A(net80),
    .VSS(VGND));
 sg13g2_inv_1 _14059_ (.VDD(VPWR),
    .Y(_00610_),
    .A(net79),
    .VSS(VGND));
 sg13g2_inv_1 _14060_ (.VDD(VPWR),
    .Y(_00611_),
    .A(net80),
    .VSS(VGND));
 sg13g2_inv_1 _14061_ (.VDD(VPWR),
    .Y(_00612_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14062_ (.VDD(VPWR),
    .Y(_00613_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14063_ (.VDD(VPWR),
    .Y(_00614_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14064_ (.VDD(VPWR),
    .Y(_00615_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14065_ (.VDD(VPWR),
    .Y(_00616_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14066_ (.VDD(VPWR),
    .Y(_00617_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14067_ (.VDD(VPWR),
    .Y(_00618_),
    .A(net95),
    .VSS(VGND));
 sg13g2_inv_1 _14068_ (.VDD(VPWR),
    .Y(_00619_),
    .A(net95),
    .VSS(VGND));
 sg13g2_inv_1 _14069_ (.VDD(VPWR),
    .Y(_00620_),
    .A(net95),
    .VSS(VGND));
 sg13g2_inv_1 _14070_ (.VDD(VPWR),
    .Y(_00621_),
    .A(net95),
    .VSS(VGND));
 sg13g2_inv_1 _14071_ (.VDD(VPWR),
    .Y(_00622_),
    .A(net95),
    .VSS(VGND));
 sg13g2_inv_1 _14072_ (.VDD(VPWR),
    .Y(_00623_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14073_ (.VDD(VPWR),
    .Y(_00624_),
    .A(net80),
    .VSS(VGND));
 sg13g2_inv_1 _14074_ (.VDD(VPWR),
    .Y(_00625_),
    .A(net94),
    .VSS(VGND));
 sg13g2_inv_1 _14075_ (.VDD(VPWR),
    .Y(_00626_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _14076_ (.VDD(VPWR),
    .Y(_00627_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _14077_ (.VDD(VPWR),
    .Y(_00628_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _14078_ (.VDD(VPWR),
    .Y(_00629_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _14079_ (.VDD(VPWR),
    .Y(_00630_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _14080_ (.VDD(VPWR),
    .Y(_00631_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _14081_ (.VDD(VPWR),
    .Y(_00632_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _14082_ (.VDD(VPWR),
    .Y(_00633_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _14083_ (.VDD(VPWR),
    .Y(_00634_),
    .A(net138),
    .VSS(VGND));
 sg13g2_inv_1 _14084_ (.VDD(VPWR),
    .Y(_00635_),
    .A(net86),
    .VSS(VGND));
 sg13g2_inv_1 _14085_ (.VDD(VPWR),
    .Y(_00636_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _14086_ (.VDD(VPWR),
    .Y(_00637_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _14087_ (.VDD(VPWR),
    .Y(_00638_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _14088_ (.VDD(VPWR),
    .Y(_00639_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14089_ (.VDD(VPWR),
    .Y(_00640_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14090_ (.VDD(VPWR),
    .Y(_00641_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14091_ (.VDD(VPWR),
    .Y(_00642_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14092_ (.VDD(VPWR),
    .Y(_00643_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14093_ (.VDD(VPWR),
    .Y(_00644_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14094_ (.VDD(VPWR),
    .Y(_00645_),
    .A(net41),
    .VSS(VGND));
 sg13g2_inv_1 _14095_ (.VDD(VPWR),
    .Y(_00646_),
    .A(net40),
    .VSS(VGND));
 sg13g2_inv_1 _14096_ (.VDD(VPWR),
    .Y(_00647_),
    .A(net41),
    .VSS(VGND));
 sg13g2_inv_1 _14097_ (.VDD(VPWR),
    .Y(_00648_),
    .A(net41),
    .VSS(VGND));
 sg13g2_inv_1 _14098_ (.VDD(VPWR),
    .Y(_00649_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _14099_ (.VDD(VPWR),
    .Y(_00650_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14100_ (.VDD(VPWR),
    .Y(_00651_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14101_ (.VDD(VPWR),
    .Y(_00652_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14102_ (.VDD(VPWR),
    .Y(_00653_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _14103_ (.VDD(VPWR),
    .Y(_00654_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14104_ (.VDD(VPWR),
    .Y(_00655_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _14105_ (.VDD(VPWR),
    .Y(_00656_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14106_ (.VDD(VPWR),
    .Y(_00657_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14107_ (.VDD(VPWR),
    .Y(_00658_),
    .A(net42),
    .VSS(VGND));
 sg13g2_inv_1 _14108_ (.VDD(VPWR),
    .Y(_00659_),
    .A(net47),
    .VSS(VGND));
 sg13g2_inv_1 _14109_ (.VDD(VPWR),
    .Y(_00660_),
    .A(net46),
    .VSS(VGND));
 sg13g2_inv_1 _14110_ (.VDD(VPWR),
    .Y(_00661_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _14111_ (.VDD(VPWR),
    .Y(_00662_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _14112_ (.VDD(VPWR),
    .Y(_00663_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _14113_ (.VDD(VPWR),
    .Y(_00664_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _14114_ (.VDD(VPWR),
    .Y(_00665_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _14115_ (.VDD(VPWR),
    .Y(_00666_),
    .A(net52),
    .VSS(VGND));
 sg13g2_inv_1 _14116_ (.VDD(VPWR),
    .Y(_00667_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _14117_ (.VDD(VPWR),
    .Y(_00668_),
    .A(net44),
    .VSS(VGND));
 sg13g2_inv_1 _14118_ (.VDD(VPWR),
    .Y(_00669_),
    .A(net46),
    .VSS(VGND));
 sg13g2_inv_1 _14119_ (.VDD(VPWR),
    .Y(_00670_),
    .A(net43),
    .VSS(VGND));
 sg13g2_inv_1 _14120_ (.VDD(VPWR),
    .Y(_00671_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _14121_ (.VDD(VPWR),
    .Y(_00672_),
    .A(net99),
    .VSS(VGND));
 sg13g2_inv_1 _14122_ (.VDD(VPWR),
    .Y(_00673_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14123_ (.VDD(VPWR),
    .Y(_00674_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14124_ (.VDD(VPWR),
    .Y(_00675_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _14125_ (.VDD(VPWR),
    .Y(_00676_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _14126_ (.VDD(VPWR),
    .Y(_00677_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _14127_ (.VDD(VPWR),
    .Y(_00678_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _14128_ (.VDD(VPWR),
    .Y(_00679_),
    .A(net119),
    .VSS(VGND));
 sg13g2_inv_1 _14129_ (.VDD(VPWR),
    .Y(_00680_),
    .A(net117),
    .VSS(VGND));
 sg13g2_inv_1 _14130_ (.VDD(VPWR),
    .Y(_00681_),
    .A(net119),
    .VSS(VGND));
 sg13g2_inv_1 _14131_ (.VDD(VPWR),
    .Y(_00682_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14132_ (.VDD(VPWR),
    .Y(_00683_),
    .A(net102),
    .VSS(VGND));
 sg13g2_inv_1 _14133_ (.VDD(VPWR),
    .Y(_00684_),
    .A(net102),
    .VSS(VGND));
 sg13g2_inv_1 _14134_ (.VDD(VPWR),
    .Y(_00685_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _14135_ (.VDD(VPWR),
    .Y(_00686_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _14136_ (.VDD(VPWR),
    .Y(_00687_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _14137_ (.VDD(VPWR),
    .Y(_00688_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _14138_ (.VDD(VPWR),
    .Y(_00689_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _14139_ (.VDD(VPWR),
    .Y(_00690_),
    .A(net89),
    .VSS(VGND));
 sg13g2_inv_1 _14140_ (.VDD(VPWR),
    .Y(_00691_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14141_ (.VDD(VPWR),
    .Y(_00692_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14142_ (.VDD(VPWR),
    .Y(_00693_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14143_ (.VDD(VPWR),
    .Y(_00694_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _14144_ (.VDD(VPWR),
    .Y(_00695_),
    .A(net129),
    .VSS(VGND));
 sg13g2_inv_1 _14145_ (.VDD(VPWR),
    .Y(_00696_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14146_ (.VDD(VPWR),
    .Y(_00697_),
    .A(net130),
    .VSS(VGND));
 sg13g2_inv_1 _14147_ (.VDD(VPWR),
    .Y(_00698_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14148_ (.VDD(VPWR),
    .Y(_00699_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14149_ (.VDD(VPWR),
    .Y(_00700_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14150_ (.VDD(VPWR),
    .Y(_00701_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14151_ (.VDD(VPWR),
    .Y(_00702_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14152_ (.VDD(VPWR),
    .Y(_00703_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14153_ (.VDD(VPWR),
    .Y(_00704_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14154_ (.VDD(VPWR),
    .Y(_00705_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14155_ (.VDD(VPWR),
    .Y(_00706_),
    .A(net130),
    .VSS(VGND));
 sg13g2_inv_1 _14156_ (.VDD(VPWR),
    .Y(_00707_),
    .A(net130),
    .VSS(VGND));
 sg13g2_inv_1 _14157_ (.VDD(VPWR),
    .Y(_00708_),
    .A(net130),
    .VSS(VGND));
 sg13g2_inv_1 _14158_ (.VDD(VPWR),
    .Y(_00709_),
    .A(net134),
    .VSS(VGND));
 sg13g2_inv_1 _14159_ (.VDD(VPWR),
    .Y(_00710_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14160_ (.VDD(VPWR),
    .Y(_00711_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14161_ (.VDD(VPWR),
    .Y(_00712_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14162_ (.VDD(VPWR),
    .Y(_00713_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14163_ (.VDD(VPWR),
    .Y(_00714_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _14164_ (.VDD(VPWR),
    .Y(_00715_),
    .A(net102),
    .VSS(VGND));
 sg13g2_inv_1 _14165_ (.VDD(VPWR),
    .Y(_00716_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14166_ (.VDD(VPWR),
    .Y(_00717_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _14167_ (.VDD(VPWR),
    .Y(_00718_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _14168_ (.VDD(VPWR),
    .Y(_00719_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14169_ (.VDD(VPWR),
    .Y(_00720_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _14170_ (.VDD(VPWR),
    .Y(_00721_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14171_ (.VDD(VPWR),
    .Y(_00722_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14172_ (.VDD(VPWR),
    .Y(_00723_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14173_ (.VDD(VPWR),
    .Y(_00724_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14174_ (.VDD(VPWR),
    .Y(_00725_),
    .A(net137),
    .VSS(VGND));
 sg13g2_inv_1 _14175_ (.VDD(VPWR),
    .Y(_00726_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _14176_ (.VDD(VPWR),
    .Y(_00727_),
    .A(net124),
    .VSS(VGND));
 sg13g2_inv_1 _14177_ (.VDD(VPWR),
    .Y(_00728_),
    .A(net127),
    .VSS(VGND));
 sg13g2_inv_1 _14178_ (.VDD(VPWR),
    .Y(_00729_),
    .A(net127),
    .VSS(VGND));
 sg13g2_inv_1 _14179_ (.VDD(VPWR),
    .Y(_00730_),
    .A(net127),
    .VSS(VGND));
 sg13g2_inv_1 _14180_ (.VDD(VPWR),
    .Y(_00731_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _14181_ (.VDD(VPWR),
    .Y(_00732_),
    .A(net139),
    .VSS(VGND));
 sg13g2_inv_1 _14182_ (.VDD(VPWR),
    .Y(_00733_),
    .A(net116),
    .VSS(VGND));
 sg13g2_inv_1 _14183_ (.VDD(VPWR),
    .Y(_00734_),
    .A(net131),
    .VSS(VGND));
 sg13g2_inv_1 _14184_ (.VDD(VPWR),
    .Y(_00735_),
    .A(net116),
    .VSS(VGND));
 sg13g2_inv_1 _14185_ (.VDD(VPWR),
    .Y(_00736_),
    .A(net116),
    .VSS(VGND));
 sg13g2_inv_1 _14186_ (.VDD(VPWR),
    .Y(_00737_),
    .A(net116),
    .VSS(VGND));
 sg13g2_inv_1 _14187_ (.VDD(VPWR),
    .Y(_00738_),
    .A(net115),
    .VSS(VGND));
 sg13g2_inv_1 _14188_ (.VDD(VPWR),
    .Y(_00739_),
    .A(net116),
    .VSS(VGND));
 sg13g2_inv_1 _14189_ (.VDD(VPWR),
    .Y(_00740_),
    .A(net104),
    .VSS(VGND));
 sg13g2_inv_1 _14190_ (.VDD(VPWR),
    .Y(_00741_),
    .A(net101),
    .VSS(VGND));
 sg13g2_inv_1 _14191_ (.VDD(VPWR),
    .Y(_00742_),
    .A(net102),
    .VSS(VGND));
 sg13g2_inv_1 _14192_ (.VDD(VPWR),
    .Y(_00743_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _14193_ (.VDD(VPWR),
    .Y(_00744_),
    .A(net91),
    .VSS(VGND));
 sg13g2_inv_1 _14194_ (.VDD(VPWR),
    .Y(_00745_),
    .A(net91),
    .VSS(VGND));
 sg13g2_inv_1 _14195_ (.VDD(VPWR),
    .Y(_00746_),
    .A(net114),
    .VSS(VGND));
 sg13g2_inv_1 _14196_ (.VDD(VPWR),
    .Y(_00747_),
    .A(net91),
    .VSS(VGND));
 sg13g2_inv_1 _14197_ (.VDD(VPWR),
    .Y(_00748_),
    .A(net90),
    .VSS(VGND));
 sg13g2_inv_1 _14198_ (.VDD(VPWR),
    .Y(_00749_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14199_ (.VDD(VPWR),
    .Y(_00750_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14200_ (.VDD(VPWR),
    .Y(_00751_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14201_ (.VDD(VPWR),
    .Y(_00752_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14202_ (.VDD(VPWR),
    .Y(_00753_),
    .A(net104),
    .VSS(VGND));
 sg13g2_inv_1 _14203_ (.VDD(VPWR),
    .Y(_00754_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14204_ (.VDD(VPWR),
    .Y(_00755_),
    .A(net103),
    .VSS(VGND));
 sg13g2_inv_1 _14205_ (.VDD(VPWR),
    .Y(_00756_),
    .A(net99),
    .VSS(VGND));
 sg13g2_inv_1 _14206_ (.VDD(VPWR),
    .Y(_00757_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14207_ (.VDD(VPWR),
    .Y(_00758_),
    .A(net106),
    .VSS(VGND));
 sg13g2_inv_1 _14208_ (.VDD(VPWR),
    .Y(_00759_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14209_ (.VDD(VPWR),
    .Y(_00760_),
    .A(net133),
    .VSS(VGND));
 sg13g2_inv_1 _14210_ (.VDD(VPWR),
    .Y(_00761_),
    .A(net135),
    .VSS(VGND));
 sg13g2_inv_1 _14211_ (.VDD(VPWR),
    .Y(_00762_),
    .A(net135),
    .VSS(VGND));
 sg13g2_inv_1 _14212_ (.VDD(VPWR),
    .Y(_00763_),
    .A(net135),
    .VSS(VGND));
 sg13g2_inv_1 _14213_ (.VDD(VPWR),
    .Y(_00764_),
    .A(net135),
    .VSS(VGND));
 sg13g2_inv_1 _14214_ (.VDD(VPWR),
    .Y(_00765_),
    .A(net133),
    .VSS(VGND));
 sg13g2_inv_1 _14215_ (.VDD(VPWR),
    .Y(_00766_),
    .A(net133),
    .VSS(VGND));
 sg13g2_inv_1 _14216_ (.VDD(VPWR),
    .Y(_00767_),
    .A(net132),
    .VSS(VGND));
 sg13g2_inv_1 _14217_ (.VDD(VPWR),
    .Y(_00768_),
    .A(net133),
    .VSS(VGND));
 sg13g2_inv_1 _14218_ (.VDD(VPWR),
    .Y(_00769_),
    .A(net105),
    .VSS(VGND));
 sg13g2_inv_1 _14219_ (.VDD(VPWR),
    .Y(_00770_),
    .A(net105),
    .VSS(VGND));
 sg13g2_dfrbpq_1 _14220_ (.RESET_B(_00021_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00771_),
    .Q(\sipo.shift_reg[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _14221_ (.RESET_B(_00022_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00772_),
    .Q(\sipo.shift_reg[2] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _14222_ (.RESET_B(_00023_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00773_),
    .Q(\sipo.shift_reg[3] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _14223_ (.RESET_B(_00024_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00774_),
    .Q(\sipo.shift_reg[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _14224_ (.RESET_B(_00025_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00775_),
    .Q(\sipo.shift_reg[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _14225_ (.RESET_B(_00026_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00776_),
    .Q(\sipo.shift_reg[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _14226_ (.RESET_B(_00027_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00777_),
    .Q(\sipo.shift_reg[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _14227_ (.RESET_B(_00028_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00778_),
    .Q(\sipo.shift_reg[8] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _14228_ (.RESET_B(_00029_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00779_),
    .Q(\sipo.shift_reg[9] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _14229_ (.RESET_B(_00030_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00780_),
    .Q(\sipo.shift_reg[10] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _14230_ (.RESET_B(_00031_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00781_),
    .Q(\sipo.shift_reg[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _14231_ (.RESET_B(_00032_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00782_),
    .Q(\sipo.shift_reg[12] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _14232_ (.RESET_B(_00033_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00783_),
    .Q(\sipo.shift_reg[13] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _14233_ (.RESET_B(_00034_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00784_),
    .Q(\sipo.shift_reg[14] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _14234_ (.RESET_B(_00035_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00785_),
    .Q(\sipo.shift_reg[15] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _14235_ (.RESET_B(_00036_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00786_),
    .Q(\instr[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14236_ (.RESET_B(_00037_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00787_),
    .Q(\instr[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _14237_ (.RESET_B(_00038_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00788_),
    .Q(\instr[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _14238_ (.RESET_B(_00039_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00789_),
    .Q(\instr[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _14239_ (.RESET_B(_00040_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00790_),
    .Q(\instr[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _14240_ (.RESET_B(_00041_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00791_),
    .Q(\instr[5] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _14241_ (.RESET_B(_00042_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00792_),
    .Q(\instr[6] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _14242_ (.RESET_B(_00043_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00793_),
    .Q(\instr[7] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _14243_ (.RESET_B(_00044_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00794_),
    .Q(\instr[8] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _14244_ (.RESET_B(_00045_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00795_),
    .Q(\instr[9] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _14245_ (.RESET_B(_00046_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00796_),
    .Q(\instr[10] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _14246_ (.RESET_B(_00047_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00797_),
    .Q(\instr[11] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _14247_ (.RESET_B(_00048_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00798_),
    .Q(\instr[12] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _14248_ (.RESET_B(_00049_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00799_),
    .Q(\instr[13] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _14249_ (.RESET_B(_00050_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00800_),
    .Q(\instr[14] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _14250_ (.RESET_B(_00051_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00801_),
    .Q(\instr[15] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _14251_ (.RESET_B(_00052_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00802_),
    .Q(\acc_sub.x2[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14252_ (.RESET_B(_00053_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00803_),
    .Q(\acc_sub.x2[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _14253_ (.RESET_B(_00054_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00804_),
    .Q(\acc_sub.x2[2] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14254_ (.RESET_B(_00055_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00805_),
    .Q(\acc_sub.x2[3] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14255_ (.RESET_B(_00056_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00806_),
    .Q(\acc_sub.x2[4] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _14256_ (.RESET_B(_00057_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00807_),
    .Q(\acc_sub.x2[5] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _14257_ (.RESET_B(_00058_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00808_),
    .Q(\acc_sub.x2[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _14258_ (.RESET_B(_00059_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00809_),
    .Q(\acc_sub.x2[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _14259_ (.RESET_B(_00060_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00810_),
    .Q(\acc_sub.x2[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _14260_ (.RESET_B(_00061_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00811_),
    .Q(\acc_sub.x2[9] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14261_ (.RESET_B(_00062_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00812_),
    .Q(\acc_sub.x2[10] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14262_ (.RESET_B(_00063_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00813_),
    .Q(\acc_sub.x2[11] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _14263_ (.RESET_B(_00064_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00814_),
    .Q(\acc_sub.x2[12] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14264_ (.RESET_B(_00065_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00815_),
    .Q(\acc_sub.x2[13] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14265_ (.RESET_B(_00066_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00816_),
    .Q(\acc_sub.x2[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _14266_ (.RESET_B(_00067_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00817_),
    .Q(\acc_sub.x2[15] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _14267_ (.RESET_B(_00068_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00818_),
    .Q(\fp16_res_pipe.x2[0] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14268_ (.RESET_B(_00069_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00819_),
    .Q(\fp16_res_pipe.x2[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _14269_ (.RESET_B(_00070_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00820_),
    .Q(\fp16_res_pipe.x2[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14270_ (.RESET_B(_00071_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00821_),
    .Q(\fp16_res_pipe.x2[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _14271_ (.RESET_B(_00072_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00822_),
    .Q(\fp16_res_pipe.x2[4] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _14272_ (.RESET_B(_00073_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00823_),
    .Q(\fp16_res_pipe.x2[5] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14273_ (.RESET_B(_00074_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00824_),
    .Q(\fp16_res_pipe.x2[6] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _14274_ (.RESET_B(_00075_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00825_),
    .Q(\fp16_res_pipe.x2[7] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14275_ (.RESET_B(_00076_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00826_),
    .Q(\fp16_res_pipe.x2[8] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _14276_ (.RESET_B(_00077_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00827_),
    .Q(\fp16_res_pipe.x2[9] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _14277_ (.RESET_B(_00078_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00828_),
    .Q(\fp16_res_pipe.x2[10] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _14278_ (.RESET_B(_00079_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00829_),
    .Q(\fp16_res_pipe.x2[11] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _14279_ (.RESET_B(_00080_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00830_),
    .Q(\fp16_res_pipe.x2[12] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _14280_ (.RESET_B(_00081_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00831_),
    .Q(\fp16_res_pipe.x2[13] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _14281_ (.RESET_B(_00082_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00832_),
    .Q(\fp16_res_pipe.x2[14] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _14282_ (.RESET_B(_00083_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00833_),
    .Q(\fp16_res_pipe.x2[15] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _14283_ (.RESET_B(_00084_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_07116_),
    .Q(\fpmul.reg1en.d[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _14284_ (.RESET_B(_00085_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_07115_),
    .Q(\fpdiv.reg1en.d[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _14285_ (.RESET_B(_00086_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_07114_),
    .Q(\fp16_sum_pipe.reg1en.d[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _14286_ (.RESET_B(_00087_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_07113_),
    .Q(\fp16_res_pipe.reg1en.d[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _14287_ (.RESET_B(_00088_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00002_),
    .Q(load_en),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _14288_ (.RESET_B(_00089_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00001_),
    .Q(\acc_sum.reg1en.d[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _14289_ (.RESET_B(_00090_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00000_),
    .Q(\acc_sub.reg1en.d[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _14290_ (.RESET_B(_00091_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00834_),
    .Q(\acc[0] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _14291_ (.RESET_B(_00092_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00835_),
    .Q(\acc[1] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _14292_ (.RESET_B(_00093_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00836_),
    .Q(\acc[2] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _14293_ (.RESET_B(_00094_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00837_),
    .Q(\acc[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _14294_ (.RESET_B(_00095_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00838_),
    .Q(\acc[4] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_2 _14295_ (.RESET_B(_00096_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00839_),
    .Q(\acc[5] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14296_ (.RESET_B(_00097_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00840_),
    .Q(\acc[6] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _14297_ (.RESET_B(_00098_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00841_),
    .Q(\acc[7] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14298_ (.RESET_B(_00099_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00842_),
    .Q(\acc[8] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14299_ (.RESET_B(_00100_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00843_),
    .Q(\acc[9] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _14300_ (.RESET_B(_00101_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00844_),
    .Q(\acc[10] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_2 _14301_ (.RESET_B(_00102_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00845_),
    .Q(\acc[11] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _14302_ (.RESET_B(_00103_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00846_),
    .Q(\acc[12] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14303_ (.RESET_B(_00104_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00847_),
    .Q(\acc[13] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _14304_ (.RESET_B(_00105_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00848_),
    .Q(\acc[14] ),
    .CLK(clknet_leaf_49_clk));
 sg13g2_dfrbpq_2 _14305_ (.RESET_B(_00106_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00849_),
    .Q(\acc[15] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _14306_ (.RESET_B(_00107_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00850_),
    .Q(\sipo.bit_counter[0] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _14307_ (.RESET_B(_00108_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00851_),
    .Q(\sipo.bit_counter[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _14308_ (.RESET_B(_00109_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00852_),
    .Q(\sipo.bit_counter[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _14309_ (.RESET_B(_00110_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00853_),
    .Q(\sipo.bit_counter[3] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _14310_ (.RESET_B(_00111_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00854_),
    .Q(\sipo.bit_counter[4] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _14311_ (.RESET_B(_00112_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00004_),
    .Q(\sipo.word_ready ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _14312_ (.RESET_B(_00113_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00855_),
    .Q(\sipo.word[0] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _14313_ (.RESET_B(_00114_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00856_),
    .Q(\sipo.word[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _14314_ (.RESET_B(_00115_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00857_),
    .Q(\sipo.word[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _14315_ (.RESET_B(_00116_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00858_),
    .Q(\sipo.word[3] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _14316_ (.RESET_B(_00117_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00859_),
    .Q(\sipo.word[4] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _14317_ (.RESET_B(_00118_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00860_),
    .Q(\sipo.word[5] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _14318_ (.RESET_B(_00119_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00861_),
    .Q(\sipo.word[6] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _14319_ (.RESET_B(_00120_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00862_),
    .Q(\sipo.word[7] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _14320_ (.RESET_B(_00121_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00863_),
    .Q(\sipo.word[8] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _14321_ (.RESET_B(_00122_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00864_),
    .Q(\sipo.word[9] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _14322_ (.RESET_B(_00123_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00865_),
    .Q(\sipo.word[10] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _14323_ (.RESET_B(_00124_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00866_),
    .Q(\sipo.word[11] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _14324_ (.RESET_B(_00125_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00867_),
    .Q(\sipo.word[12] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _14325_ (.RESET_B(_00126_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00868_),
    .Q(\sipo.word[13] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _14326_ (.RESET_B(_00127_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00869_),
    .Q(\sipo.word[14] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _14327_ (.RESET_B(_00128_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00870_),
    .Q(\sipo.word[15] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _14328_ (.RESET_B(_00129_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00871_),
    .Q(\piso.tx_active ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _14329_ (.RESET_B(_00130_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00003_),
    .Q(\sipo.receiving ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _14330_ (.RESET_B(_00131_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00872_),
    .Q(net4),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _14331_ (.RESET_B(_00132_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00873_),
    .Q(\piso.tx_bit_counter[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _14332_ (.RESET_B(_00133_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00874_),
    .Q(\piso.tx_bit_counter[1] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _14333_ (.RESET_B(_00134_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00875_),
    .Q(\piso.tx_bit_counter[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _14334_ (.RESET_B(_00135_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00876_),
    .Q(\piso.tx_bit_counter[3] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _14335_ (.RESET_B(_00136_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00877_),
    .Q(\piso.tx_bit_counter[4] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_1 _14336_ (.RESET_B(_00137_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00878_),
    .Q(\fpmul.reg_p_out[0] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _14337_ (.RESET_B(_00138_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00879_),
    .Q(\fpmul.reg_p_out[1] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _14338_ (.RESET_B(_00139_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00880_),
    .Q(\fpmul.reg_p_out[2] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _14339_ (.RESET_B(_00140_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00881_),
    .Q(\fpmul.reg_p_out[3] ),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _14340_ (.RESET_B(_00141_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00882_),
    .Q(\fpmul.reg_p_out[4] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _14341_ (.RESET_B(_00142_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00883_),
    .Q(\fpmul.reg_p_out[5] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _14342_ (.RESET_B(_00143_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00884_),
    .Q(\fpmul.reg_p_out[6] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _14343_ (.RESET_B(_00144_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00885_),
    .Q(\fpmul.reg_p_out[7] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _14344_ (.RESET_B(_00145_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00886_),
    .Q(\fpmul.reg_p_out[8] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _14345_ (.RESET_B(_00146_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00887_),
    .Q(\fpmul.reg_p_out[9] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _14346_ (.RESET_B(_00147_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00888_),
    .Q(\fpmul.reg_p_out[10] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _14347_ (.RESET_B(_00148_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00889_),
    .Q(\fpmul.reg_p_out[11] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _14348_ (.RESET_B(_00149_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00890_),
    .Q(\fpmul.reg_p_out[12] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _14349_ (.RESET_B(_00150_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00891_),
    .Q(\fpmul.reg_p_out[13] ),
    .CLK(clknet_leaf_94_clk));
 sg13g2_dfrbpq_1 _14350_ (.RESET_B(_00151_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00892_),
    .Q(\fpmul.reg_p_out[14] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _14351_ (.RESET_B(_00152_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00893_),
    .Q(\fpmul.reg_p_out[15] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _14352_ (.RESET_B(_00153_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00894_),
    .Q(_00005_),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _14353_ (.RESET_B(_00154_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00895_),
    .Q(_00006_),
    .CLK(clknet_leaf_82_clk));
 sg13g2_dfrbpq_1 _14354_ (.RESET_B(_00155_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00896_),
    .Q(_00007_),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14355_ (.RESET_B(_00156_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00897_),
    .Q(_00008_),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14356_ (.RESET_B(_00157_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00898_),
    .Q(_00009_),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14357_ (.RESET_B(_00158_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00899_),
    .Q(_00010_),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _14358_ (.RESET_B(_00159_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00900_),
    .Q(_00011_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14359_ (.RESET_B(_00160_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00901_),
    .Q(_00012_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14360_ (.RESET_B(_00161_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00902_),
    .Q(_00013_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14361_ (.RESET_B(_00162_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00903_),
    .Q(_00014_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14362_ (.RESET_B(_00163_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00904_),
    .Q(_00015_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14363_ (.RESET_B(_00164_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00905_),
    .Q(_00016_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14364_ (.RESET_B(_00165_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00906_),
    .Q(_00017_),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _14365_ (.RESET_B(_00166_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00907_),
    .Q(_00018_),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14366_ (.RESET_B(_00167_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00908_),
    .Q(_00019_),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _14367_ (.RESET_B(_00168_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00909_),
    .Q(_00020_),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_2 _14368_ (.RESET_B(_00169_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1955),
    .Q(\fpmul.reg1en.q[0] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _14369_ (.RESET_B(_00170_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00910_),
    .Q(\fpmul.reg_b_out[0] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_2 _14370_ (.RESET_B(_00171_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00911_),
    .Q(\fpmul.reg_b_out[1] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_1 _14371_ (.RESET_B(_00172_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00912_),
    .Q(\fpmul.reg_b_out[2] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _14372_ (.RESET_B(_00173_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00913_),
    .Q(\fpmul.reg_b_out[3] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _14373_ (.RESET_B(_00174_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00914_),
    .Q(\fpmul.reg_b_out[4] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _14374_ (.RESET_B(_00175_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00915_),
    .Q(\fpmul.reg_b_out[5] ),
    .CLK(clknet_leaf_106_clk));
 sg13g2_dfrbpq_2 _14375_ (.RESET_B(_00176_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00916_),
    .Q(\fpmul.reg_b_out[6] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_2 _14376_ (.RESET_B(_00177_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00917_),
    .Q(\fpmul.reg_b_out[7] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _14377_ (.RESET_B(_00178_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00918_),
    .Q(\fpmul.reg_b_out[8] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _14378_ (.RESET_B(_00179_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00919_),
    .Q(\fpmul.reg_b_out[9] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _14379_ (.RESET_B(_00180_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00920_),
    .Q(\fpmul.reg_b_out[10] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _14380_ (.RESET_B(_00181_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00921_),
    .Q(\fpmul.reg_b_out[11] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _14381_ (.RESET_B(_00182_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00922_),
    .Q(\fpmul.reg_b_out[12] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _14382_ (.RESET_B(_00183_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00923_),
    .Q(\fpmul.reg_b_out[13] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _14383_ (.RESET_B(_00184_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00924_),
    .Q(\fpmul.reg_b_out[14] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_1 _14384_ (.RESET_B(_00185_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00925_),
    .Q(\fpmul.reg_b_out[15] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _14385_ (.RESET_B(_00186_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1873),
    .Q(\fpmul.reg2en.q[0] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _14386_ (.RESET_B(_00187_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1861),
    .Q(\fpmul.reg3en.q[0] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _14387_ (.RESET_B(_00188_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00926_),
    .Q(\div_result[0] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _14388_ (.RESET_B(_00189_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00927_),
    .Q(\div_result[1] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _14389_ (.RESET_B(_00190_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00928_),
    .Q(\div_result[2] ),
    .CLK(clknet_leaf_83_clk));
 sg13g2_dfrbpq_1 _14390_ (.RESET_B(_00191_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00929_),
    .Q(\div_result[3] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14391_ (.RESET_B(_00192_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00930_),
    .Q(\div_result[4] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _14392_ (.RESET_B(_00193_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00931_),
    .Q(\div_result[5] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_1 _14393_ (.RESET_B(_00194_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00932_),
    .Q(\div_result[6] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14394_ (.RESET_B(_00195_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00933_),
    .Q(\div_result[7] ),
    .CLK(clknet_leaf_88_clk));
 sg13g2_dfrbpq_1 _14395_ (.RESET_B(_00196_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00934_),
    .Q(\div_result[8] ),
    .CLK(clknet_leaf_87_clk));
 sg13g2_dfrbpq_1 _14396_ (.RESET_B(_00197_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00935_),
    .Q(\div_result[9] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _14397_ (.RESET_B(_00198_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00936_),
    .Q(\div_result[10] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _14398_ (.RESET_B(_00199_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00937_),
    .Q(\div_result[11] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _14399_ (.RESET_B(_00200_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00938_),
    .Q(\div_result[12] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _14400_ (.RESET_B(_00201_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00939_),
    .Q(\div_result[13] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _14401_ (.RESET_B(_00202_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00940_),
    .Q(\div_result[14] ),
    .CLK(clknet_leaf_89_clk));
 sg13g2_dfrbpq_1 _14402_ (.RESET_B(_00203_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00941_),
    .Q(\div_result[15] ),
    .CLK(clknet_leaf_90_clk));
 sg13g2_dfrbpq_1 _14403_ (.RESET_B(_00204_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00942_),
    .Q(\fpmul.reg_a_out[0] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _14404_ (.RESET_B(_00205_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00943_),
    .Q(\fpmul.reg_a_out[1] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _14405_ (.RESET_B(_00206_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00944_),
    .Q(\fpmul.reg_a_out[2] ),
    .CLK(clknet_leaf_102_clk));
 sg13g2_dfrbpq_2 _14406_ (.RESET_B(_00207_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00945_),
    .Q(\fpmul.reg_a_out[3] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _14407_ (.RESET_B(_00208_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00946_),
    .Q(\fpmul.reg_a_out[4] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _14408_ (.RESET_B(_00209_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00947_),
    .Q(\fpmul.reg_a_out[5] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _14409_ (.RESET_B(_00210_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00948_),
    .Q(\fpmul.reg_a_out[6] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_2 _14410_ (.RESET_B(_00211_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00949_),
    .Q(\fpmul.reg_a_out[7] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14411_ (.RESET_B(_00212_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00950_),
    .Q(\fpmul.reg_a_out[8] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _14412_ (.RESET_B(_00213_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00951_),
    .Q(\fpmul.reg_a_out[9] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_2 _14413_ (.RESET_B(_00214_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00952_),
    .Q(\fpmul.reg_a_out[10] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14414_ (.RESET_B(_00215_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00953_),
    .Q(\fpmul.reg_a_out[11] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _14415_ (.RESET_B(_00216_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00954_),
    .Q(\fpmul.reg_a_out[12] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14416_ (.RESET_B(_00217_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00955_),
    .Q(\fpmul.reg_a_out[13] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_2 _14417_ (.RESET_B(_00218_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00956_),
    .Q(\fpmul.reg_a_out[14] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _14418_ (.RESET_B(_00219_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00957_),
    .Q(\fpmul.reg_a_out[15] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_1 _14419_ (.RESET_B(_00220_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00958_),
    .Q(\fpmul.seg_reg0.q[4] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _14420_ (.RESET_B(_00221_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00959_),
    .Q(\fpmul.seg_reg0.q[5] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _14421_ (.RESET_B(_00222_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00960_),
    .Q(\fpmul.seg_reg0.q[6] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _14422_ (.RESET_B(_00223_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00961_),
    .Q(\fpmul.seg_reg0.q[7] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _14423_ (.RESET_B(_00224_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00962_),
    .Q(\fpmul.seg_reg0.q[8] ),
    .CLK(clknet_leaf_79_clk));
 sg13g2_dfrbpq_1 _14424_ (.RESET_B(_00225_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00963_),
    .Q(\fpmul.seg_reg0.q[9] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _14425_ (.RESET_B(_00226_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00964_),
    .Q(\fpmul.seg_reg0.q[10] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _14426_ (.RESET_B(_00227_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00965_),
    .Q(\fpmul.seg_reg0.q[11] ),
    .CLK(clknet_leaf_78_clk));
 sg13g2_dfrbpq_1 _14427_ (.RESET_B(_00228_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00966_),
    .Q(\fpmul.seg_reg0.q[12] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _14428_ (.RESET_B(_00229_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00967_),
    .Q(\fpmul.seg_reg0.q[13] ),
    .CLK(clknet_leaf_80_clk));
 sg13g2_dfrbpq_1 _14429_ (.RESET_B(_00230_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00968_),
    .Q(\fpmul.seg_reg0.q[14] ),
    .CLK(clknet_leaf_81_clk));
 sg13g2_dfrbpq_2 _14430_ (.RESET_B(_00231_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00969_),
    .Q(\fpmul.seg_reg0.q[15] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _14431_ (.RESET_B(_00232_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00970_),
    .Q(\fpmul.seg_reg0.q[16] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _14432_ (.RESET_B(_00233_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00971_),
    .Q(\fpmul.seg_reg0.q[17] ),
    .CLK(clknet_leaf_101_clk));
 sg13g2_dfrbpq_1 _14433_ (.RESET_B(_00234_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00972_),
    .Q(\fpmul.seg_reg0.q[18] ),
    .CLK(clknet_leaf_95_clk));
 sg13g2_dfrbpq_1 _14434_ (.RESET_B(_00235_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00973_),
    .Q(\fpmul.seg_reg0.q[19] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _14435_ (.RESET_B(_00236_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00974_),
    .Q(\fpmul.seg_reg0.q[20] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _14436_ (.RESET_B(_00237_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00975_),
    .Q(\fpmul.seg_reg0.q[21] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _14437_ (.RESET_B(_00238_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00976_),
    .Q(\fpmul.seg_reg0.q[22] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _14438_ (.RESET_B(_00239_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00977_),
    .Q(\fpmul.seg_reg0.q[23] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _14439_ (.RESET_B(_00240_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00978_),
    .Q(\fpmul.seg_reg0.q[24] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _14440_ (.RESET_B(_00241_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00979_),
    .Q(\fpmul.seg_reg0.q[25] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _14441_ (.RESET_B(_00242_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00980_),
    .Q(\fpmul.seg_reg0.q[26] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _14442_ (.RESET_B(_00243_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00981_),
    .Q(\fpmul.seg_reg0.q[27] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _14443_ (.RESET_B(_00244_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00982_),
    .Q(\fpmul.seg_reg0.q[28] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _14444_ (.RESET_B(_00245_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00983_),
    .Q(\fpmul.seg_reg0.q[29] ),
    .CLK(clknet_leaf_105_clk));
 sg13g2_dfrbpq_1 _14445_ (.RESET_B(_00246_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00984_),
    .Q(\fpmul.seg_reg0.q[30] ),
    .CLK(clknet_leaf_103_clk));
 sg13g2_dfrbpq_1 _14446_ (.RESET_B(_00247_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00985_),
    .Q(\fpmul.seg_reg0.q[31] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _14447_ (.RESET_B(_00248_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00986_),
    .Q(\fpmul.seg_reg0.q[32] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _14448_ (.RESET_B(_00249_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00987_),
    .Q(\fpmul.seg_reg0.q[33] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _14449_ (.RESET_B(_00250_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00988_),
    .Q(\fpmul.seg_reg0.q[34] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_1 _14450_ (.RESET_B(_00251_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00989_),
    .Q(\fpmul.seg_reg0.q[35] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _14451_ (.RESET_B(_00252_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00990_),
    .Q(\fpmul.seg_reg0.q[36] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _14452_ (.RESET_B(_00253_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00991_),
    .Q(\fpmul.seg_reg0.q[37] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _14453_ (.RESET_B(_00254_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00992_),
    .Q(\fpmul.seg_reg0.q[38] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _14454_ (.RESET_B(_00255_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00993_),
    .Q(\fpmul.seg_reg0.q[39] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _14455_ (.RESET_B(_00256_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00994_),
    .Q(\fpmul.seg_reg0.q[40] ),
    .CLK(clknet_leaf_104_clk));
 sg13g2_dfrbpq_1 _14456_ (.RESET_B(_00257_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00995_),
    .Q(\fpmul.seg_reg0.q[41] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _14457_ (.RESET_B(_00258_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00996_),
    .Q(\fpmul.seg_reg0.q[42] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _14458_ (.RESET_B(_00259_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00997_),
    .Q(\fpmul.seg_reg0.q[43] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _14459_ (.RESET_B(_00260_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00998_),
    .Q(\fpmul.seg_reg0.q[44] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _14460_ (.RESET_B(_00261_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_00999_),
    .Q(\fpmul.seg_reg0.q[45] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _14461_ (.RESET_B(_00262_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01000_),
    .Q(\fpmul.seg_reg0.q[46] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _14462_ (.RESET_B(_00263_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01001_),
    .Q(\fpmul.seg_reg0.q[47] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _14463_ (.RESET_B(_00264_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01002_),
    .Q(\fpmul.seg_reg0.q[48] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _14464_ (.RESET_B(_00265_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01003_),
    .Q(\fpmul.seg_reg0.q[49] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _14465_ (.RESET_B(_00266_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01004_),
    .Q(\fpmul.seg_reg0.q[50] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_1 _14466_ (.RESET_B(_00267_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01005_),
    .Q(\fpmul.seg_reg0.q[51] ),
    .CLK(clknet_leaf_93_clk));
 sg13g2_dfrbpq_1 _14467_ (.RESET_B(_00268_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01006_),
    .Q(\fpmul.seg_reg0.q[52] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _14468_ (.RESET_B(_00269_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01007_),
    .Q(\fpmul.seg_reg0.q[53] ),
    .CLK(clknet_leaf_125_clk));
 sg13g2_dfrbpq_1 _14469_ (.RESET_B(_00270_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01008_),
    .Q(\fpmul.result[15] ),
    .CLK(clknet_leaf_92_clk));
 sg13g2_dfrbpq_1 _14470_ (.RESET_B(_00271_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01009_),
    .Q(\fpdiv.divider0.counter[0] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_1 _14471_ (.RESET_B(_00272_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01010_),
    .Q(\fpdiv.divider0.counter[1] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _14472_ (.RESET_B(_00273_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01011_),
    .Q(\fpdiv.divider0.counter[2] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _14473_ (.RESET_B(_00274_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01012_),
    .Q(\fpdiv.divider0.counter[3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _14474_ (.RESET_B(_00275_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\fpdiv.divider0.en_r ),
    .Q(\fpdiv.divider0.state ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _14475_ (.RESET_B(_00276_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01013_),
    .Q(\add_result[0] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _14476_ (.RESET_B(_00277_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01014_),
    .Q(\add_result[1] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_1 _14477_ (.RESET_B(_00278_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01015_),
    .Q(\add_result[2] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _14478_ (.RESET_B(_00279_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01016_),
    .Q(\add_result[3] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _14479_ (.RESET_B(_00280_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01017_),
    .Q(\add_result[4] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _14480_ (.RESET_B(_00281_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01018_),
    .Q(\add_result[5] ),
    .CLK(clknet_leaf_107_clk));
 sg13g2_dfrbpq_1 _14481_ (.RESET_B(_00282_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01019_),
    .Q(\add_result[6] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_1 _14482_ (.RESET_B(_00283_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01020_),
    .Q(\add_result[7] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _14483_ (.RESET_B(_00284_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01021_),
    .Q(\add_result[8] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _14484_ (.RESET_B(_00285_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01022_),
    .Q(\add_result[9] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _14485_ (.RESET_B(_00286_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01023_),
    .Q(\add_result[10] ),
    .CLK(clknet_leaf_100_clk));
 sg13g2_dfrbpq_2 _14486_ (.RESET_B(_00287_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01024_),
    .Q(\add_result[11] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _14487_ (.RESET_B(_00288_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01025_),
    .Q(\add_result[12] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _14488_ (.RESET_B(_00289_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01026_),
    .Q(\add_result[13] ),
    .CLK(clknet_leaf_99_clk));
 sg13g2_dfrbpq_2 _14489_ (.RESET_B(_00290_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01027_),
    .Q(\add_result[14] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _14490_ (.RESET_B(_00291_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01028_),
    .Q(\add_result[15] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14491_ (.RESET_B(_00292_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1741),
    .Q(\fpdiv.reg2en.q[0] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _14492_ (.RESET_B(_00293_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1947),
    .Q(\fpdiv.reg1en.q[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_2 _14493_ (.RESET_B(_00294_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01029_),
    .Q(\fpdiv.divider0.divisor[4] ),
    .CLK(clknet_leaf_86_clk));
 sg13g2_dfrbpq_1 _14494_ (.RESET_B(_00295_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01030_),
    .Q(\fpdiv.divider0.divisor[5] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _14495_ (.RESET_B(_00296_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01031_),
    .Q(\fpdiv.divider0.divisor[6] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _14496_ (.RESET_B(_00297_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01032_),
    .Q(\fpdiv.divider0.divisor[7] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14497_ (.RESET_B(_00298_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01033_),
    .Q(\fpdiv.divider0.divisor[8] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _14498_ (.RESET_B(_00299_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01034_),
    .Q(\fpdiv.divider0.divisor[9] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_1 _14499_ (.RESET_B(_00300_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01035_),
    .Q(\fpdiv.divider0.divisor[10] ),
    .CLK(clknet_leaf_84_clk));
 sg13g2_dfrbpq_2 _14500_ (.RESET_B(_00301_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01036_),
    .Q(\fpdiv.reg_b_out[7] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _14501_ (.RESET_B(_00302_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01037_),
    .Q(\fpdiv.reg_b_out[8] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _14502_ (.RESET_B(_00303_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01038_),
    .Q(\fpdiv.reg_b_out[9] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _14503_ (.RESET_B(_00304_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01039_),
    .Q(\fpdiv.reg_b_out[10] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _14504_ (.RESET_B(_00305_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01040_),
    .Q(\fpdiv.reg_b_out[11] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _14505_ (.RESET_B(_00306_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01041_),
    .Q(\fpdiv.reg_b_out[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _14506_ (.RESET_B(_00307_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01042_),
    .Q(\fpdiv.reg_b_out[13] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _14507_ (.RESET_B(_00308_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01043_),
    .Q(\fpdiv.reg_b_out[14] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _14508_ (.RESET_B(_00309_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01044_),
    .Q(\fpdiv.reg_b_out[15] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _14509_ (.RESET_B(_00310_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01045_),
    .Q(\fpdiv.divider0.dividend[4] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _14510_ (.RESET_B(_00311_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01046_),
    .Q(\fpdiv.divider0.dividend[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _14511_ (.RESET_B(_00312_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01047_),
    .Q(\fpdiv.divider0.dividend[6] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_1 _14512_ (.RESET_B(_00313_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01048_),
    .Q(\fpdiv.divider0.dividend[7] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _14513_ (.RESET_B(_00314_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01049_),
    .Q(\fpdiv.divider0.dividend[8] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_1 _14514_ (.RESET_B(_00315_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01050_),
    .Q(\fpdiv.divider0.dividend[9] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _14515_ (.RESET_B(_00316_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01051_),
    .Q(\fpdiv.divider0.dividend[10] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _14516_ (.RESET_B(_00317_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01052_),
    .Q(\fpdiv.reg_a_out[7] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _14517_ (.RESET_B(_00318_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01053_),
    .Q(\fpdiv.reg_a_out[8] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_2 _14518_ (.RESET_B(_00319_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01054_),
    .Q(\fpdiv.reg_a_out[9] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _14519_ (.RESET_B(_00320_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01055_),
    .Q(\fpdiv.reg_a_out[10] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _14520_ (.RESET_B(_00321_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01056_),
    .Q(\fpdiv.reg_a_out[11] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_1 _14521_ (.RESET_B(_00322_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01057_),
    .Q(\fpdiv.reg_a_out[12] ),
    .CLK(clknet_leaf_53_clk));
 sg13g2_dfrbpq_2 _14522_ (.RESET_B(_00323_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01058_),
    .Q(\fpdiv.reg_a_out[13] ),
    .CLK(clknet_leaf_126_clk));
 sg13g2_dfrbpq_2 _14523_ (.RESET_B(_00324_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01059_),
    .Q(\fpdiv.reg_a_out[14] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _14524_ (.RESET_B(_00325_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01060_),
    .Q(\fpdiv.reg_a_out[15] ),
    .CLK(clknet_leaf_91_clk));
 sg13g2_dfrbpq_1 _14525_ (.RESET_B(_00326_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01061_),
    .Q(\fpdiv.div_out[0] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _14526_ (.RESET_B(_00327_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01062_),
    .Q(\fpdiv.div_out[1] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _14527_ (.RESET_B(_00328_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01063_),
    .Q(\fpdiv.div_out[2] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_1 _14528_ (.RESET_B(_00329_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01064_),
    .Q(\fpdiv.div_out[3] ),
    .CLK(clknet_leaf_72_clk));
 sg13g2_dfrbpq_2 _14529_ (.RESET_B(_00330_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01065_),
    .Q(\fpdiv.div_out[4] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _14530_ (.RESET_B(_00331_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01066_),
    .Q(\fpdiv.div_out[5] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _14531_ (.RESET_B(_00332_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01067_),
    .Q(\fpdiv.div_out[6] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _14532_ (.RESET_B(_00333_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01068_),
    .Q(\fpdiv.div_out[7] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _14533_ (.RESET_B(_00334_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01069_),
    .Q(\fpdiv.div_out[8] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_1 _14534_ (.RESET_B(_00335_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01070_),
    .Q(\fpdiv.div_out[9] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_1 _14535_ (.RESET_B(_00336_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01071_),
    .Q(\fpdiv.div_out[10] ),
    .CLK(clknet_leaf_76_clk));
 sg13g2_dfrbpq_2 _14536_ (.RESET_B(_00337_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01072_),
    .Q(\fpdiv.div_out[11] ),
    .CLK(clknet_leaf_77_clk));
 sg13g2_dfrbpq_2 _14537_ (.RESET_B(_00338_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01073_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _14538_ (.RESET_B(_00339_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01074_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[1] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _14539_ (.RESET_B(_00340_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01075_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _14540_ (.RESET_B(_00341_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01076_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _14541_ (.RESET_B(_00342_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01077_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _14542_ (.RESET_B(_00343_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01078_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _14543_ (.RESET_B(_00344_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01079_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[6] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _14544_ (.RESET_B(_00345_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01080_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[7] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _14545_ (.RESET_B(_00346_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01081_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[8] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _14546_ (.RESET_B(_00347_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01082_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[9] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _14547_ (.RESET_B(_00348_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01083_),
    .Q(\acc_sum.op_sign_logic0.mantisa_b[10] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _14548_ (.RESET_B(_00349_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01084_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[0] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _14549_ (.RESET_B(_00350_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01085_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[1] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _14550_ (.RESET_B(_00351_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01086_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[2] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _14551_ (.RESET_B(_00352_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01087_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[3] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _14552_ (.RESET_B(_00353_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01088_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[4] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _14553_ (.RESET_B(_00354_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01089_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[5] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _14554_ (.RESET_B(_00355_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01090_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[6] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _14555_ (.RESET_B(_00356_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01091_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[7] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_2 _14556_ (.RESET_B(_00357_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01092_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[8] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _14557_ (.RESET_B(_00358_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01093_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[9] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _14558_ (.RESET_B(_00359_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01094_),
    .Q(\acc_sum.op_sign_logic0.mantisa_a[10] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _14559_ (.RESET_B(_00360_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01095_),
    .Q(\acc_sum.seg_reg0.q[22] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _14560_ (.RESET_B(_00361_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01096_),
    .Q(\acc_sum.seg_reg0.q[23] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _14561_ (.RESET_B(_00362_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01097_),
    .Q(\acc_sum.seg_reg0.q[24] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _14562_ (.RESET_B(_00363_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01098_),
    .Q(\acc_sum.seg_reg0.q[25] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _14563_ (.RESET_B(_00364_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01099_),
    .Q(\acc_sum.seg_reg0.q[26] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_2 _14564_ (.RESET_B(_00365_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01100_),
    .Q(\acc_sum.seg_reg0.q[27] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _14565_ (.RESET_B(_00366_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01101_),
    .Q(\acc_sum.seg_reg0.q[28] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _14566_ (.RESET_B(_00367_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01102_),
    .Q(\acc_sum.seg_reg0.q[29] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _14567_ (.RESET_B(_00368_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01103_),
    .Q(\acc_sum.op_sign_logic0.s_b ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _14568_ (.RESET_B(_00369_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01104_),
    .Q(\acc_sum.op_sign_logic0.s_a ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _14569_ (.RESET_B(_00370_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\fp16_sum_pipe.reg3en.q[0] ),
    .Q(\fp16_sum_pipe.reg4en.q[0] ),
    .CLK(clknet_leaf_96_clk));
 sg13g2_dfrbpq_2 _14570_ (.RESET_B(_00371_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1846),
    .Q(\fp16_sum_pipe.reg3en.q[0] ),
    .CLK(clknet_leaf_97_clk));
 sg13g2_dfrbpq_2 _14571_ (.RESET_B(_00372_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1843),
    .Q(\fp16_sum_pipe.reg2en.q[0] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _14572_ (.RESET_B(_00373_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1933),
    .Q(\fp16_sum_pipe.reg1en.q[0] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _14573_ (.RESET_B(_00374_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01105_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[0] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _14574_ (.RESET_B(_00375_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01106_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[1] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _14575_ (.RESET_B(_00376_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01107_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[2] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _14576_ (.RESET_B(_00377_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01108_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[3] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_2 _14577_ (.RESET_B(_00378_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01109_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[4] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_1 _14578_ (.RESET_B(_00379_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01110_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[5] ),
    .CLK(clknet_leaf_117_clk));
 sg13g2_dfrbpq_2 _14579_ (.RESET_B(_00380_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01111_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[6] ),
    .CLK(clknet_leaf_135_clk));
 sg13g2_dfrbpq_1 _14580_ (.RESET_B(_00381_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01112_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[7] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _14581_ (.RESET_B(_00382_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01113_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[8] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _14582_ (.RESET_B(_00383_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01114_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[9] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14583_ (.RESET_B(_00384_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01115_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[10] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_1 _14584_ (.RESET_B(_00385_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01116_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[11] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _14585_ (.RESET_B(_00386_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01117_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[12] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _14586_ (.RESET_B(_00387_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01118_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[13] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _14587_ (.RESET_B(_00388_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01119_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[14] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_1 _14588_ (.RESET_B(_00389_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01120_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.b[15] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14589_ (.RESET_B(_00390_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01121_),
    .Q(\fp16_res_pipe.y[0] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _14590_ (.RESET_B(_00391_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01122_),
    .Q(\fp16_res_pipe.y[1] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_1 _14591_ (.RESET_B(_00392_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01123_),
    .Q(\fp16_res_pipe.y[2] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _14592_ (.RESET_B(_00393_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01124_),
    .Q(\fp16_res_pipe.y[3] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _14593_ (.RESET_B(_00394_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01125_),
    .Q(\fp16_res_pipe.y[4] ),
    .CLK(clknet_leaf_127_clk));
 sg13g2_dfrbpq_2 _14594_ (.RESET_B(_00395_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01126_),
    .Q(\fp16_res_pipe.y[5] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _14595_ (.RESET_B(_00396_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01127_),
    .Q(\fp16_res_pipe.y[6] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _14596_ (.RESET_B(_00397_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01128_),
    .Q(\fp16_res_pipe.y[7] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _14597_ (.RESET_B(_00398_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01129_),
    .Q(\fp16_res_pipe.y[8] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_1 _14598_ (.RESET_B(_00399_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01130_),
    .Q(\fp16_res_pipe.y[9] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _14599_ (.RESET_B(_00400_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01131_),
    .Q(\fp16_res_pipe.y[10] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _14600_ (.RESET_B(_00401_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01132_),
    .Q(\fp16_res_pipe.y[11] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _14601_ (.RESET_B(_00402_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01133_),
    .Q(\fp16_res_pipe.y[12] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _14602_ (.RESET_B(_00403_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01134_),
    .Q(\fp16_res_pipe.y[13] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_1 _14603_ (.RESET_B(_00404_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01135_),
    .Q(\fp16_res_pipe.y[14] ),
    .CLK(clknet_leaf_129_clk));
 sg13g2_dfrbpq_2 _14604_ (.RESET_B(_00405_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01136_),
    .Q(\fp16_res_pipe.y[15] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _14605_ (.RESET_B(_00406_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01137_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[0] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _14606_ (.RESET_B(_00407_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01138_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[1] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _14607_ (.RESET_B(_00408_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01139_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[2] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _14608_ (.RESET_B(_00409_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01140_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[3] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _14609_ (.RESET_B(_00410_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01141_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[4] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _14610_ (.RESET_B(_00411_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01142_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[5] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_2 _14611_ (.RESET_B(_00412_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01143_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[6] ),
    .CLK(clknet_leaf_118_clk));
 sg13g2_dfrbpq_2 _14612_ (.RESET_B(_00413_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01144_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[7] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _14613_ (.RESET_B(_00414_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01145_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[8] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _14614_ (.RESET_B(_00415_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01146_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[9] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14615_ (.RESET_B(_00416_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01147_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[10] ),
    .CLK(clknet_leaf_122_clk));
 sg13g2_dfrbpq_2 _14616_ (.RESET_B(_00417_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01148_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[11] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _14617_ (.RESET_B(_00418_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01149_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[12] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_1 _14618_ (.RESET_B(_00419_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01150_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[13] ),
    .CLK(clknet_leaf_123_clk));
 sg13g2_dfrbpq_2 _14619_ (.RESET_B(_00420_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01151_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[14] ),
    .CLK(clknet_leaf_134_clk));
 sg13g2_dfrbpq_2 _14620_ (.RESET_B(_00421_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01152_),
    .Q(\fp16_sum_pipe.exp_mant_logic0.a[15] ),
    .CLK(clknet_leaf_124_clk));
 sg13g2_dfrbpq_2 _14621_ (.RESET_B(_00422_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01153_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[0] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_2 _14622_ (.RESET_B(_00423_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01154_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[1] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _14623_ (.RESET_B(_00424_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01155_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[2] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _14624_ (.RESET_B(_00425_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01156_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[3] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _14625_ (.RESET_B(_00426_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01157_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[4] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_1 _14626_ (.RESET_B(_00427_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01158_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[5] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_2 _14627_ (.RESET_B(_00428_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01159_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[6] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _14628_ (.RESET_B(_00429_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01160_),
    .Q(\fp16_sum_pipe.add_renorm0.exp[7] ),
    .CLK(clknet_leaf_98_clk));
 sg13g2_dfrbpq_1 _14629_ (.RESET_B(_00430_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01161_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[0] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _14630_ (.RESET_B(_00431_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01162_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[1] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _14631_ (.RESET_B(_00432_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01163_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[2] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _14632_ (.RESET_B(_00433_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01164_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[3] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _14633_ (.RESET_B(_00434_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01165_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[4] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _14634_ (.RESET_B(_00435_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01166_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[5] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _14635_ (.RESET_B(_00436_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01167_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[6] ),
    .CLK(clknet_leaf_108_clk));
 sg13g2_dfrbpq_2 _14636_ (.RESET_B(_00437_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01168_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[7] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_1 _14637_ (.RESET_B(_00438_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01169_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[8] ),
    .CLK(clknet_leaf_109_clk));
 sg13g2_dfrbpq_2 _14638_ (.RESET_B(_00439_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01170_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[9] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _14639_ (.RESET_B(_00440_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01171_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[10] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_2 _14640_ (.RESET_B(_00441_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01172_),
    .Q(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .CLK(clknet_leaf_110_clk));
 sg13g2_dfrbpq_1 _14641_ (.RESET_B(_00442_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01173_),
    .Q(\fp16_sum_pipe.seg_reg1.q[20] ),
    .CLK(clknet_leaf_120_clk));
 sg13g2_dfrbpq_2 _14642_ (.RESET_B(_00443_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01174_),
    .Q(\fp16_sum_pipe.seg_reg1.q[21] ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _14643_ (.RESET_B(_00444_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1835),
    .Q(\fp16_res_pipe.reg4en.q[0] ),
    .CLK(clknet_leaf_128_clk));
 sg13g2_dfrbpq_2 _14644_ (.RESET_B(_00445_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1833),
    .Q(\fp16_res_pipe.reg3en.q[0] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _14645_ (.RESET_B(_00446_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\fp16_res_pipe.reg1en.q[0] ),
    .Q(\fp16_res_pipe.reg2en.q[0] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _14646_ (.RESET_B(_00447_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1916),
    .Q(\fp16_res_pipe.reg1en.q[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _14647_ (.RESET_B(_00448_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01175_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[0] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _14648_ (.RESET_B(_00449_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01176_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _14649_ (.RESET_B(_00450_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01177_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[2] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _14650_ (.RESET_B(_00451_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01178_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[3] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _14651_ (.RESET_B(_00452_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01179_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[4] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_2 _14652_ (.RESET_B(_00453_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01180_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[5] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _14653_ (.RESET_B(_00454_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01181_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[6] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_1 _14654_ (.RESET_B(_00455_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01182_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[7] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _14655_ (.RESET_B(_00456_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01183_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[8] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _14656_ (.RESET_B(_00457_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01184_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[9] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _14657_ (.RESET_B(_00458_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01185_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[10] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _14658_ (.RESET_B(_00459_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01186_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _14659_ (.RESET_B(_00460_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01187_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _14660_ (.RESET_B(_00461_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01188_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[13] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _14661_ (.RESET_B(_00462_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01189_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[14] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _14662_ (.RESET_B(_00463_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01190_),
    .Q(\fp16_res_pipe.exp_mant_logic0.b[15] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _14663_ (.RESET_B(_00464_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01191_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[0] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _14664_ (.RESET_B(_00465_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01192_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[1] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _14665_ (.RESET_B(_00466_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01193_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[2] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _14666_ (.RESET_B(_00467_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01194_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[3] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _14667_ (.RESET_B(_00468_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01195_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[4] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_2 _14668_ (.RESET_B(_00469_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01196_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[5] ),
    .CLK(clknet_leaf_141_clk));
 sg13g2_dfrbpq_2 _14669_ (.RESET_B(_00470_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01197_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[6] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _14670_ (.RESET_B(_00471_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01198_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[7] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _14671_ (.RESET_B(_00472_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01199_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[8] ),
    .CLK(clknet_leaf_140_clk));
 sg13g2_dfrbpq_1 _14672_ (.RESET_B(_00473_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01200_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[9] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _14673_ (.RESET_B(_00474_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01201_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_b[10] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _14674_ (.RESET_B(_00475_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01202_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[0] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _14675_ (.RESET_B(_00476_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01203_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[1] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _14676_ (.RESET_B(_00477_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01204_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[2] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _14677_ (.RESET_B(_00478_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01205_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _14678_ (.RESET_B(_00479_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01206_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[4] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _14679_ (.RESET_B(_00480_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01207_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[5] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _14680_ (.RESET_B(_00481_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01208_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[6] ),
    .CLK(clknet_leaf_144_clk));
 sg13g2_dfrbpq_2 _14681_ (.RESET_B(_00482_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01209_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[7] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _14682_ (.RESET_B(_00483_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01210_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[8] ),
    .CLK(clknet_leaf_143_clk));
 sg13g2_dfrbpq_2 _14683_ (.RESET_B(_00484_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01211_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[9] ),
    .CLK(clknet_leaf_142_clk));
 sg13g2_dfrbpq_1 _14684_ (.RESET_B(_00485_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01212_),
    .Q(\fp16_res_pipe.op_sign_logic0.mantisa_a[10] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _14685_ (.RESET_B(_00486_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01213_),
    .Q(\fp16_res_pipe.seg_reg0.q[22] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _14686_ (.RESET_B(_00487_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01214_),
    .Q(\fp16_res_pipe.seg_reg0.q[23] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _14687_ (.RESET_B(_00488_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01215_),
    .Q(\fp16_res_pipe.seg_reg0.q[24] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _14688_ (.RESET_B(_00489_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01216_),
    .Q(\fp16_res_pipe.seg_reg0.q[25] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _14689_ (.RESET_B(_00490_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01217_),
    .Q(\fp16_res_pipe.seg_reg0.q[26] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _14690_ (.RESET_B(_00491_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01218_),
    .Q(\fp16_res_pipe.seg_reg0.q[27] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _14691_ (.RESET_B(_00492_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01219_),
    .Q(\fp16_res_pipe.seg_reg0.q[28] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _14692_ (.RESET_B(_00493_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01220_),
    .Q(\fp16_res_pipe.seg_reg0.q[29] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _14693_ (.RESET_B(_00494_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01221_),
    .Q(\fp16_res_pipe.op_sign_logic0.add_sub ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _14694_ (.RESET_B(_00495_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01222_),
    .Q(\fp16_res_pipe.op_sign_logic0.s_b ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _14695_ (.RESET_B(_00496_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01223_),
    .Q(\fp16_res_pipe.op_sign_logic0.s_a ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _14696_ (.RESET_B(_00497_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01224_),
    .Q(\fp16_res_pipe.reg_add_sub.q[0] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_1 _14697_ (.RESET_B(_00498_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01225_),
    .Q(\acc_sum.y[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _14698_ (.RESET_B(_00499_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01226_),
    .Q(\acc_sum.y[1] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _14699_ (.RESET_B(_00500_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01227_),
    .Q(\acc_sum.y[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _14700_ (.RESET_B(_00501_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01228_),
    .Q(\acc_sum.y[3] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _14701_ (.RESET_B(_00502_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01229_),
    .Q(\acc_sum.y[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _14702_ (.RESET_B(_00503_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01230_),
    .Q(\acc_sum.y[5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _14703_ (.RESET_B(_00504_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01231_),
    .Q(\acc_sum.y[6] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _14704_ (.RESET_B(_00505_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01232_),
    .Q(\acc_sum.y[7] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _14705_ (.RESET_B(_00506_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01233_),
    .Q(\acc_sum.y[8] ),
    .CLK(clknet_leaf_47_clk));
 sg13g2_dfrbpq_1 _14706_ (.RESET_B(_00507_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01234_),
    .Q(\acc_sum.y[9] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _14707_ (.RESET_B(_00508_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01235_),
    .Q(\acc_sum.y[10] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _14708_ (.RESET_B(_00509_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01236_),
    .Q(\acc_sum.y[11] ),
    .CLK(clknet_leaf_48_clk));
 sg13g2_dfrbpq_1 _14709_ (.RESET_B(_00510_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01237_),
    .Q(\acc_sum.y[12] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _14710_ (.RESET_B(_00511_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01238_),
    .Q(\acc_sum.y[13] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _14711_ (.RESET_B(_00512_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01239_),
    .Q(\acc_sum.y[14] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _14712_ (.RESET_B(_00513_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01240_),
    .Q(\acc_sum.y[15] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _14713_ (.RESET_B(_00514_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01241_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _14714_ (.RESET_B(_00515_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01242_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _14715_ (.RESET_B(_00516_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01243_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[2] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _14716_ (.RESET_B(_00517_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01244_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _14717_ (.RESET_B(_00518_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01245_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _14718_ (.RESET_B(_00519_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01246_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _14719_ (.RESET_B(_00520_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01247_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _14720_ (.RESET_B(_00521_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01248_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[7] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _14721_ (.RESET_B(_00522_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01249_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[8] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _14722_ (.RESET_B(_00523_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01250_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[9] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_2 _14723_ (.RESET_B(_00524_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01251_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[10] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _14724_ (.RESET_B(_00525_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01252_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[11] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _14725_ (.RESET_B(_00526_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01253_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[12] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _14726_ (.RESET_B(_00527_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01254_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[13] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _14727_ (.RESET_B(_00528_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01255_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[14] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _14728_ (.RESET_B(_00529_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01256_),
    .Q(\fp16_res_pipe.exp_mant_logic0.a[15] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _14729_ (.RESET_B(_00530_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01257_),
    .Q(\fp16_res_pipe.add_renorm0.exp[0] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _14730_ (.RESET_B(_00531_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01258_),
    .Q(\fp16_res_pipe.add_renorm0.exp[1] ),
    .CLK(clknet_5_2__leaf_clk));
 sg13g2_dfrbpq_1 _14731_ (.RESET_B(_00532_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01259_),
    .Q(\fp16_res_pipe.add_renorm0.exp[2] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _14732_ (.RESET_B(_00533_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01260_),
    .Q(\fp16_res_pipe.add_renorm0.exp[3] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_1 _14733_ (.RESET_B(_00534_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01261_),
    .Q(\fp16_res_pipe.add_renorm0.exp[4] ),
    .CLK(clknet_leaf_132_clk));
 sg13g2_dfrbpq_2 _14734_ (.RESET_B(_00535_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01262_),
    .Q(\fp16_res_pipe.add_renorm0.exp[5] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _14735_ (.RESET_B(_00536_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01263_),
    .Q(\fp16_res_pipe.add_renorm0.exp[6] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _14736_ (.RESET_B(_00537_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01264_),
    .Q(\fp16_res_pipe.add_renorm0.exp[7] ),
    .CLK(clknet_leaf_131_clk));
 sg13g2_dfrbpq_1 _14737_ (.RESET_B(_00538_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01265_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[0] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _14738_ (.RESET_B(_00539_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01266_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[1] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _14739_ (.RESET_B(_00540_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01267_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[2] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _14740_ (.RESET_B(_00541_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01268_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[3] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _14741_ (.RESET_B(_00542_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01269_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[4] ),
    .CLK(clknet_5_0__leaf_clk));
 sg13g2_dfrbpq_2 _14742_ (.RESET_B(_00543_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01270_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[5] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _14743_ (.RESET_B(_00544_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01271_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[6] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_2 _14744_ (.RESET_B(_00545_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01272_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[7] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _14745_ (.RESET_B(_00546_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01273_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[8] ),
    .CLK(clknet_leaf_136_clk));
 sg13g2_dfrbpq_2 _14746_ (.RESET_B(_00547_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01274_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[9] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _14747_ (.RESET_B(_00548_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01275_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[10] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_2 _14748_ (.RESET_B(_00549_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01276_),
    .Q(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .CLK(clknet_leaf_137_clk));
 sg13g2_dfrbpq_1 _14749_ (.RESET_B(_00550_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01277_),
    .Q(\fp16_res_pipe.seg_reg1.q[20] ),
    .CLK(clknet_leaf_130_clk));
 sg13g2_dfrbpq_2 _14750_ (.RESET_B(_00551_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01278_),
    .Q(\fp16_res_pipe.seg_reg1.q[21] ),
    .CLK(clknet_leaf_139_clk));
 sg13g2_dfrbpq_1 _14751_ (.RESET_B(_00552_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(\acc_sum.reg3en.q[0] ),
    .Q(\acc_sum.reg4en.q[0] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _14752_ (.RESET_B(_00553_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1819),
    .Q(\acc_sum.reg3en.q[0] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _14753_ (.RESET_B(_00554_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1813),
    .Q(\acc_sum.reg2en.q[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _14754_ (.RESET_B(_00555_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1899),
    .Q(\acc_sum.reg1en.q[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _14755_ (.RESET_B(_00556_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01279_),
    .Q(\acc_sum.exp_mant_logic0.b[0] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _14756_ (.RESET_B(_00557_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01280_),
    .Q(\acc_sum.exp_mant_logic0.b[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _14757_ (.RESET_B(_00558_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01281_),
    .Q(\acc_sum.exp_mant_logic0.b[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _14758_ (.RESET_B(_00559_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01282_),
    .Q(\acc_sum.exp_mant_logic0.b[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _14759_ (.RESET_B(_00560_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01283_),
    .Q(\acc_sum.exp_mant_logic0.b[4] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _14760_ (.RESET_B(_00561_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01284_),
    .Q(\acc_sum.exp_mant_logic0.b[5] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _14761_ (.RESET_B(_00562_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01285_),
    .Q(\acc_sum.exp_mant_logic0.b[6] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _14762_ (.RESET_B(_00563_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01286_),
    .Q(\acc_sum.exp_mant_logic0.b[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _14763_ (.RESET_B(_00564_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01287_),
    .Q(\acc_sum.exp_mant_logic0.b[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _14764_ (.RESET_B(_00565_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01288_),
    .Q(\acc_sum.exp_mant_logic0.b[9] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _14765_ (.RESET_B(_00566_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01289_),
    .Q(\acc_sum.exp_mant_logic0.b[10] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _14766_ (.RESET_B(_00567_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01290_),
    .Q(\acc_sum.exp_mant_logic0.b[11] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _14767_ (.RESET_B(_00568_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01291_),
    .Q(\acc_sum.exp_mant_logic0.b[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _14768_ (.RESET_B(_00569_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01292_),
    .Q(\acc_sum.exp_mant_logic0.b[13] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _14769_ (.RESET_B(_00570_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01293_),
    .Q(\acc_sum.exp_mant_logic0.b[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _14770_ (.RESET_B(_00571_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01294_),
    .Q(\acc_sum.exp_mant_logic0.b[15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _14771_ (.RESET_B(_00572_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01295_),
    .Q(\acc_sub.y[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _14772_ (.RESET_B(_00573_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01296_),
    .Q(\acc_sub.y[1] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14773_ (.RESET_B(_00574_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01297_),
    .Q(\acc_sub.y[2] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14774_ (.RESET_B(_00575_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01298_),
    .Q(\acc_sub.y[3] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14775_ (.RESET_B(_00576_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01299_),
    .Q(\acc_sub.y[4] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14776_ (.RESET_B(_00577_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01300_),
    .Q(\acc_sub.y[5] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _14777_ (.RESET_B(_00578_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01301_),
    .Q(\acc_sub.y[6] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14778_ (.RESET_B(_00579_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01302_),
    .Q(\acc_sub.y[7] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14779_ (.RESET_B(_00580_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01303_),
    .Q(\acc_sub.y[8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _14780_ (.RESET_B(_00581_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01304_),
    .Q(\acc_sub.y[9] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _14781_ (.RESET_B(_00582_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01305_),
    .Q(\acc_sub.y[10] ),
    .CLK(clknet_5_21__leaf_clk));
 sg13g2_dfrbpq_1 _14782_ (.RESET_B(_00583_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01306_),
    .Q(\acc_sub.y[11] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _14783_ (.RESET_B(_00584_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01307_),
    .Q(\acc_sub.y[12] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _14784_ (.RESET_B(_00585_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01308_),
    .Q(\acc_sub.y[13] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _14785_ (.RESET_B(_00586_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01309_),
    .Q(\acc_sub.y[14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _14786_ (.RESET_B(_00587_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01310_),
    .Q(\acc_sub.y[15] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_2 _14787_ (.RESET_B(_00588_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01311_),
    .Q(\acc_sum.exp_mant_logic0.a[0] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _14788_ (.RESET_B(_00589_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01312_),
    .Q(\acc_sum.exp_mant_logic0.a[1] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _14789_ (.RESET_B(_00590_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01313_),
    .Q(\acc_sum.exp_mant_logic0.a[2] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _14790_ (.RESET_B(_00591_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01314_),
    .Q(\acc_sum.exp_mant_logic0.a[3] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _14791_ (.RESET_B(_00592_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01315_),
    .Q(\acc_sum.exp_mant_logic0.a[4] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _14792_ (.RESET_B(_00593_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01316_),
    .Q(\acc_sum.exp_mant_logic0.a[5] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _14793_ (.RESET_B(_00594_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01317_),
    .Q(\acc_sum.exp_mant_logic0.a[6] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _14794_ (.RESET_B(_00595_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01318_),
    .Q(\acc_sum.exp_mant_logic0.a[7] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_2 _14795_ (.RESET_B(_00596_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01319_),
    .Q(\acc_sum.exp_mant_logic0.a[8] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _14796_ (.RESET_B(_00597_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01320_),
    .Q(\acc_sum.exp_mant_logic0.a[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _14797_ (.RESET_B(_00598_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01321_),
    .Q(\acc_sum.exp_mant_logic0.a[10] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _14798_ (.RESET_B(_00599_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01322_),
    .Q(\acc_sum.exp_mant_logic0.a[11] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _14799_ (.RESET_B(_00600_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01323_),
    .Q(\acc_sum.exp_mant_logic0.a[12] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _14800_ (.RESET_B(_00601_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01324_),
    .Q(\acc_sum.exp_mant_logic0.a[13] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _14801_ (.RESET_B(_00602_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01325_),
    .Q(\acc_sum.exp_mant_logic0.a[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _14802_ (.RESET_B(_00603_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01326_),
    .Q(\acc_sum.exp_mant_logic0.a[15] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _14803_ (.RESET_B(_00604_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01327_),
    .Q(\acc_sum.add_renorm0.exp[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _14804_ (.RESET_B(_00605_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01328_),
    .Q(\acc_sum.add_renorm0.exp[1] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _14805_ (.RESET_B(_00606_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01329_),
    .Q(\acc_sum.add_renorm0.exp[2] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _14806_ (.RESET_B(_00607_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01330_),
    .Q(\acc_sum.add_renorm0.exp[3] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _14807_ (.RESET_B(_00608_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01331_),
    .Q(\acc_sum.add_renorm0.exp[4] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _14808_ (.RESET_B(_00609_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01332_),
    .Q(\acc_sum.add_renorm0.exp[5] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _14809_ (.RESET_B(_00610_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01333_),
    .Q(\acc_sum.add_renorm0.exp[6] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _14810_ (.RESET_B(_00611_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01334_),
    .Q(\acc_sum.add_renorm0.exp[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _14811_ (.RESET_B(_00612_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01335_),
    .Q(\acc_sum.add_renorm0.mantisa[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _14812_ (.RESET_B(_00613_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01336_),
    .Q(\acc_sum.add_renorm0.mantisa[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _14813_ (.RESET_B(_00614_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01337_),
    .Q(\acc_sum.add_renorm0.mantisa[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _14814_ (.RESET_B(_00615_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01338_),
    .Q(\acc_sum.add_renorm0.mantisa[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _14815_ (.RESET_B(_00616_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01339_),
    .Q(\acc_sum.add_renorm0.mantisa[4] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _14816_ (.RESET_B(_00617_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01340_),
    .Q(\acc_sum.add_renorm0.mantisa[5] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _14817_ (.RESET_B(_00618_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01341_),
    .Q(\acc_sum.add_renorm0.mantisa[6] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _14818_ (.RESET_B(_00619_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01342_),
    .Q(\acc_sum.add_renorm0.mantisa[7] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _14819_ (.RESET_B(_00620_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01343_),
    .Q(\acc_sum.add_renorm0.mantisa[8] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _14820_ (.RESET_B(_00621_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01344_),
    .Q(\acc_sum.add_renorm0.mantisa[9] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_2 _14821_ (.RESET_B(_00622_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01345_),
    .Q(\acc_sum.add_renorm0.mantisa[10] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _14822_ (.RESET_B(_00623_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01346_),
    .Q(\acc_sum.add_renorm0.mantisa[11] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _14823_ (.RESET_B(_00624_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01347_),
    .Q(\acc_sum.seg_reg1.q[20] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _14824_ (.RESET_B(_00625_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01348_),
    .Q(\acc_sum.seg_reg1.q[21] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _14825_ (.RESET_B(_00626_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01349_),
    .Q(\fpdiv.divider0.remainder_reg[4] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _14826_ (.RESET_B(_00627_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01350_),
    .Q(\fpdiv.divider0.remainder_reg[5] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _14827_ (.RESET_B(_00628_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01351_),
    .Q(\fpdiv.divider0.remainder_reg[6] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _14828_ (.RESET_B(_00629_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01352_),
    .Q(\fpdiv.divider0.remainder_reg[7] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_2 _14829_ (.RESET_B(_00630_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01353_),
    .Q(\fpdiv.divider0.remainder_reg[8] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _14830_ (.RESET_B(_00631_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01354_),
    .Q(\fpdiv.divider0.remainder_reg[9] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _14831_ (.RESET_B(_00632_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01355_),
    .Q(\fpdiv.divider0.remainder_reg[10] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _14832_ (.RESET_B(_00633_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01356_),
    .Q(\fpdiv.divider0.remainder_reg[11] ),
    .CLK(clknet_leaf_73_clk));
 sg13g2_dfrbpq_1 _14833_ (.RESET_B(_00634_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01357_),
    .Q(\fpdiv.divider0.remainder_reg[12] ),
    .CLK(clknet_leaf_71_clk));
 sg13g2_dfrbpq_2 _14834_ (.RESET_B(_00635_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01358_),
    .Q(\state[0] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _14835_ (.RESET_B(_00636_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01359_),
    .Q(\state[1] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_2 _14836_ (.RESET_B(_00637_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01360_),
    .Q(\state[2] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _14837_ (.RESET_B(_00638_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01361_),
    .Q(\state[3] ),
    .CLK(clknet_leaf_52_clk));
 sg13g2_dfrbpq_1 _14838_ (.RESET_B(_00639_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01362_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[0] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _14839_ (.RESET_B(_00640_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01363_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[1] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _14840_ (.RESET_B(_00641_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01364_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[2] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _14841_ (.RESET_B(_00642_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01365_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[3] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _14842_ (.RESET_B(_00643_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01366_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[4] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _14843_ (.RESET_B(_00644_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01367_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[5] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _14844_ (.RESET_B(_00645_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01368_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[6] ),
    .CLK(clknet_leaf_116_clk));
 sg13g2_dfrbpq_2 _14845_ (.RESET_B(_00646_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01369_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[7] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _14846_ (.RESET_B(_00647_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01370_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[8] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_2 _14847_ (.RESET_B(_00648_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01371_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[9] ),
    .CLK(clknet_leaf_115_clk));
 sg13g2_dfrbpq_1 _14848_ (.RESET_B(_00649_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01372_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_b[10] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _14849_ (.RESET_B(_00650_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01373_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[0] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _14850_ (.RESET_B(_00651_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01374_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[1] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_2 _14851_ (.RESET_B(_00652_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01375_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[2] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _14852_ (.RESET_B(_00653_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01376_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[3] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_2 _14853_ (.RESET_B(_00654_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01377_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[4] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _14854_ (.RESET_B(_00655_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01378_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[5] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _14855_ (.RESET_B(_00656_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01379_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[6] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _14856_ (.RESET_B(_00657_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01380_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[7] ),
    .CLK(clknet_leaf_114_clk));
 sg13g2_dfrbpq_1 _14857_ (.RESET_B(_00658_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01381_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[8] ),
    .CLK(clknet_5_8__leaf_clk));
 sg13g2_dfrbpq_1 _14858_ (.RESET_B(_00659_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01382_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[9] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _14859_ (.RESET_B(_00660_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01383_),
    .Q(\fp16_sum_pipe.op_sign_logic0.mantisa_a[10] ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _14860_ (.RESET_B(_00661_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01384_),
    .Q(\fp16_sum_pipe.seg_reg0.q[22] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14861_ (.RESET_B(_00662_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01385_),
    .Q(\fp16_sum_pipe.seg_reg0.q[23] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14862_ (.RESET_B(_00663_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01386_),
    .Q(\fp16_sum_pipe.seg_reg0.q[24] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _14863_ (.RESET_B(_00664_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01387_),
    .Q(\fp16_sum_pipe.seg_reg0.q[25] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14864_ (.RESET_B(_00665_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01388_),
    .Q(\fp16_sum_pipe.seg_reg0.q[26] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _14865_ (.RESET_B(_00666_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01389_),
    .Q(\fp16_sum_pipe.seg_reg0.q[27] ),
    .CLK(clknet_leaf_121_clk));
 sg13g2_dfrbpq_1 _14866_ (.RESET_B(_00667_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01390_),
    .Q(\fp16_sum_pipe.seg_reg0.q[28] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _14867_ (.RESET_B(_00668_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01391_),
    .Q(\fp16_sum_pipe.seg_reg0.q[29] ),
    .CLK(clknet_leaf_119_clk));
 sg13g2_dfrbpq_1 _14868_ (.RESET_B(_00669_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01392_),
    .Q(\fp16_sum_pipe.op_sign_logic0.s_b ),
    .CLK(clknet_leaf_111_clk));
 sg13g2_dfrbpq_1 _14869_ (.RESET_B(_00670_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01393_),
    .Q(\fp16_sum_pipe.op_sign_logic0.s_a ),
    .CLK(clknet_leaf_112_clk));
 sg13g2_dfrbpq_1 _14870_ (.RESET_B(_00671_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1800),
    .Q(\acc_sub.reg4en.q[0] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _14871_ (.RESET_B(_00672_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1797),
    .Q(\acc_sub.reg3en.q[0] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_2 _14872_ (.RESET_B(_00673_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1796),
    .Q(\acc_sub.reg2en.q[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _14873_ (.RESET_B(_00674_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1895),
    .Q(\acc_sub.reg1en.q[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _14874_ (.RESET_B(_00675_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01394_),
    .Q(\acc_sub.exp_mant_logic0.b[0] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _14875_ (.RESET_B(_00676_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01395_),
    .Q(\acc_sub.exp_mant_logic0.b[1] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _14876_ (.RESET_B(_00677_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01396_),
    .Q(\acc_sub.exp_mant_logic0.b[2] ),
    .CLK(clknet_leaf_57_clk));
 sg13g2_dfrbpq_2 _14877_ (.RESET_B(_00678_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01397_),
    .Q(\acc_sub.exp_mant_logic0.b[3] ),
    .CLK(clknet_leaf_59_clk));
 sg13g2_dfrbpq_2 _14878_ (.RESET_B(_00679_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01398_),
    .Q(\acc_sub.exp_mant_logic0.b[4] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _14879_ (.RESET_B(_00680_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01399_),
    .Q(\acc_sub.exp_mant_logic0.b[5] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_2 _14880_ (.RESET_B(_00681_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01400_),
    .Q(\acc_sub.exp_mant_logic0.b[6] ),
    .CLK(clknet_leaf_58_clk));
 sg13g2_dfrbpq_1 _14881_ (.RESET_B(_00682_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01401_),
    .Q(\acc_sub.exp_mant_logic0.b[7] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _14882_ (.RESET_B(_00683_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01402_),
    .Q(\acc_sub.exp_mant_logic0.b[8] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _14883_ (.RESET_B(_00684_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01403_),
    .Q(\acc_sub.exp_mant_logic0.b[9] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_2 _14884_ (.RESET_B(_00685_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01404_),
    .Q(\acc_sub.exp_mant_logic0.b[10] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _14885_ (.RESET_B(_00686_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01405_),
    .Q(\acc_sub.exp_mant_logic0.b[11] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _14886_ (.RESET_B(_00687_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01406_),
    .Q(\acc_sub.exp_mant_logic0.b[12] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_2 _14887_ (.RESET_B(_00688_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01407_),
    .Q(\acc_sub.exp_mant_logic0.b[13] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_2 _14888_ (.RESET_B(_00689_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01408_),
    .Q(\acc_sub.exp_mant_logic0.b[14] ),
    .CLK(clknet_leaf_54_clk));
 sg13g2_dfrbpq_1 _14889_ (.RESET_B(_00690_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01409_),
    .Q(\acc_sub.exp_mant_logic0.b[15] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _14890_ (.RESET_B(_00691_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01410_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _14891_ (.RESET_B(_00692_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01411_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[1] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _14892_ (.RESET_B(_00693_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01412_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[2] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _14893_ (.RESET_B(_00694_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01413_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[3] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _14894_ (.RESET_B(_00695_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01414_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[4] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_1 _14895_ (.RESET_B(_00696_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01415_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[5] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _14896_ (.RESET_B(_00697_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01416_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[6] ),
    .CLK(clknet_leaf_69_clk));
 sg13g2_dfrbpq_2 _14897_ (.RESET_B(_00698_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01417_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[7] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _14898_ (.RESET_B(_00699_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01418_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[8] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_2 _14899_ (.RESET_B(_00700_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01419_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[9] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _14900_ (.RESET_B(_00701_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01420_),
    .Q(\acc_sub.op_sign_logic0.mantisa_b[10] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _14901_ (.RESET_B(_00702_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01421_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_2 _14902_ (.RESET_B(_00703_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01422_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[1] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _14903_ (.RESET_B(_00704_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01423_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _14904_ (.RESET_B(_00705_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01424_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[3] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _14905_ (.RESET_B(_00706_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01425_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[4] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _14906_ (.RESET_B(_00707_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01426_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[5] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_2 _14907_ (.RESET_B(_00708_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01427_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[6] ),
    .CLK(clknet_leaf_68_clk));
 sg13g2_dfrbpq_1 _14908_ (.RESET_B(_00709_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01428_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[7] ),
    .CLK(clknet_leaf_67_clk));
 sg13g2_dfrbpq_1 _14909_ (.RESET_B(_00710_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01429_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[8] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _14910_ (.RESET_B(_00711_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01430_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[9] ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_1 _14911_ (.RESET_B(_00712_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01431_),
    .Q(\acc_sub.op_sign_logic0.mantisa_a[10] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _14912_ (.RESET_B(_00713_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01432_),
    .Q(\acc_sub.seg_reg0.q[22] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _14913_ (.RESET_B(_00714_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01433_),
    .Q(\acc_sub.seg_reg0.q[23] ),
    .CLK(clknet_leaf_46_clk));
 sg13g2_dfrbpq_1 _14914_ (.RESET_B(_00715_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01434_),
    .Q(\acc_sub.seg_reg0.q[24] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _14915_ (.RESET_B(_00716_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01435_),
    .Q(\acc_sub.seg_reg0.q[25] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _14916_ (.RESET_B(_00717_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01436_),
    .Q(\acc_sub.seg_reg0.q[26] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_1 _14917_ (.RESET_B(_00718_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01437_),
    .Q(\acc_sub.seg_reg0.q[27] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _14918_ (.RESET_B(_00719_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01438_),
    .Q(\acc_sub.seg_reg0.q[28] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _14919_ (.RESET_B(_00720_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01439_),
    .Q(\acc_sub.seg_reg0.q[29] ),
    .CLK(clknet_leaf_50_clk));
 sg13g2_dfrbpq_2 _14920_ (.RESET_B(_00721_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01440_),
    .Q(\acc_sub.op_sign_logic0.add_sub ),
    .CLK(clknet_leaf_62_clk));
 sg13g2_dfrbpq_2 _14921_ (.RESET_B(_00722_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01441_),
    .Q(\acc_sub.op_sign_logic0.s_b ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _14922_ (.RESET_B(_00723_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01442_),
    .Q(\acc_sub.op_sign_logic0.s_a ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _14923_ (.RESET_B(_00724_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01443_),
    .Q(\acc_sub.reg_add_sub.q[0] ),
    .CLK(clknet_leaf_61_clk));
 sg13g2_dfrbpq_1 _14924_ (.RESET_B(_00725_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01444_),
    .Q(\fpdiv.divider0.divisor_reg[4] ),
    .CLK(clknet_leaf_74_clk));
 sg13g2_dfrbpq_1 _14925_ (.RESET_B(_00726_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01445_),
    .Q(\fpdiv.divider0.divisor_reg[5] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _14926_ (.RESET_B(_00727_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01446_),
    .Q(\fpdiv.divider0.divisor_reg[6] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_2 _14927_ (.RESET_B(_00728_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01447_),
    .Q(\fpdiv.divider0.divisor_reg[7] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _14928_ (.RESET_B(_00729_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01448_),
    .Q(\fpdiv.divider0.divisor_reg[8] ),
    .CLK(clknet_leaf_85_clk));
 sg13g2_dfrbpq_2 _14929_ (.RESET_B(_00730_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01449_),
    .Q(\fpdiv.divider0.divisor_reg[9] ),
    .CLK(clknet_leaf_75_clk));
 sg13g2_dfrbpq_1 _14930_ (.RESET_B(_00731_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01450_),
    .Q(\fpdiv.divider0.divisor_reg[10] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_1 _14931_ (.RESET_B(_00732_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01451_),
    .Q(\fpdiv.divider0.divisor_reg[11] ),
    .CLK(clknet_leaf_70_clk));
 sg13g2_dfrbpq_2 _14932_ (.RESET_B(_00733_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01452_),
    .Q(\acc_sub.exp_mant_logic0.a[0] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _14933_ (.RESET_B(_00734_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01453_),
    .Q(\acc_sub.exp_mant_logic0.a[1] ),
    .CLK(clknet_5_28__leaf_clk));
 sg13g2_dfrbpq_2 _14934_ (.RESET_B(_00735_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01454_),
    .Q(\acc_sub.exp_mant_logic0.a[2] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _14935_ (.RESET_B(_00736_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01455_),
    .Q(\acc_sub.exp_mant_logic0.a[3] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _14936_ (.RESET_B(_00737_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01456_),
    .Q(\acc_sub.exp_mant_logic0.a[4] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _14937_ (.RESET_B(_00738_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01457_),
    .Q(\acc_sub.exp_mant_logic0.a[5] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_2 _14938_ (.RESET_B(_00739_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01458_),
    .Q(\acc_sub.exp_mant_logic0.a[6] ),
    .CLK(clknet_leaf_56_clk));
 sg13g2_dfrbpq_1 _14939_ (.RESET_B(_00740_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01459_),
    .Q(\acc_sub.exp_mant_logic0.a[7] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _14940_ (.RESET_B(_00741_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01460_),
    .Q(\acc_sub.exp_mant_logic0.a[8] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _14941_ (.RESET_B(_00742_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01461_),
    .Q(\acc_sub.exp_mant_logic0.a[9] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _14942_ (.RESET_B(_00743_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01462_),
    .Q(\acc_sub.exp_mant_logic0.a[10] ),
    .CLK(clknet_leaf_45_clk));
 sg13g2_dfrbpq_1 _14943_ (.RESET_B(_00744_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01463_),
    .Q(\acc_sub.exp_mant_logic0.a[11] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _14944_ (.RESET_B(_00745_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01464_),
    .Q(\acc_sub.exp_mant_logic0.a[12] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_1 _14945_ (.RESET_B(_00746_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01465_),
    .Q(\acc_sub.exp_mant_logic0.a[13] ),
    .CLK(clknet_leaf_55_clk));
 sg13g2_dfrbpq_1 _14946_ (.RESET_B(_00747_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01466_),
    .Q(\acc_sub.exp_mant_logic0.a[14] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _14947_ (.RESET_B(_00748_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01467_),
    .Q(\acc_sub.exp_mant_logic0.a[15] ),
    .CLK(clknet_leaf_51_clk));
 sg13g2_dfrbpq_2 _14948_ (.RESET_B(_00749_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01468_),
    .Q(\acc_sub.add_renorm0.exp[0] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _14949_ (.RESET_B(_00750_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01469_),
    .Q(\acc_sub.add_renorm0.exp[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _14950_ (.RESET_B(_00751_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01470_),
    .Q(\acc_sub.add_renorm0.exp[2] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _14951_ (.RESET_B(_00752_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01471_),
    .Q(\acc_sub.add_renorm0.exp[3] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _14952_ (.RESET_B(_00753_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01472_),
    .Q(\acc_sub.add_renorm0.exp[4] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _14953_ (.RESET_B(_00754_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01473_),
    .Q(\acc_sub.add_renorm0.exp[5] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _14954_ (.RESET_B(_00755_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01474_),
    .Q(\acc_sub.add_renorm0.exp[6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _14955_ (.RESET_B(_00756_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01475_),
    .Q(\acc_sub.add_renorm0.exp[7] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _14956_ (.RESET_B(_00757_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01476_),
    .Q(\acc_sub.add_renorm0.mantisa[0] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _14957_ (.RESET_B(_00758_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01477_),
    .Q(\acc_sub.add_renorm0.mantisa[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_2 _14958_ (.RESET_B(_00759_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01478_),
    .Q(\acc_sub.add_renorm0.mantisa[2] ),
    .CLK(clknet_5_29__leaf_clk));
 sg13g2_dfrbpq_2 _14959_ (.RESET_B(_00760_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01479_),
    .Q(\acc_sub.add_renorm0.mantisa[3] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _14960_ (.RESET_B(_00761_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01480_),
    .Q(\acc_sub.add_renorm0.mantisa[4] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _14961_ (.RESET_B(_00762_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01481_),
    .Q(\acc_sub.add_renorm0.mantisa[5] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _14962_ (.RESET_B(_00763_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01482_),
    .Q(\acc_sub.add_renorm0.mantisa[6] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _14963_ (.RESET_B(_00764_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01483_),
    .Q(\acc_sub.add_renorm0.mantisa[7] ),
    .CLK(clknet_leaf_66_clk));
 sg13g2_dfrbpq_2 _14964_ (.RESET_B(_00765_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01484_),
    .Q(\acc_sub.add_renorm0.mantisa[8] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _14965_ (.RESET_B(_00766_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01485_),
    .Q(\acc_sub.add_renorm0.mantisa[9] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_2 _14966_ (.RESET_B(_00767_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01486_),
    .Q(\acc_sub.add_renorm0.mantisa[10] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _14967_ (.RESET_B(_00768_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01487_),
    .Q(\acc_sub.add_renorm0.mantisa[11] ),
    .CLK(clknet_leaf_63_clk));
 sg13g2_dfrbpq_1 _14968_ (.RESET_B(_00769_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01488_),
    .Q(\acc_sub.seg_reg1.q[20] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _14969_ (.RESET_B(_00770_),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_01489_),
    .Q(\acc_sub.seg_reg1.q[21] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_buf_2 place1639 (.A(_02352_),
    .X(net1639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1640 (.A(_02063_),
    .X(net1640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1641 (.A(_01944_),
    .X(net1641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1642 (.A(_04190_),
    .X(net1642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1643 (.A(_04158_),
    .X(net1643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1644 (.A(_04126_),
    .X(net1644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1645 (.A(_02324_),
    .X(net1645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1646 (.A(_01949_),
    .X(net1646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1651 (.A(_01923_),
    .X(net1651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1652 (.A(_02322_),
    .X(net1652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1654 (.A(_05141_),
    .X(net1654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_81_clk (.A(clknet_5_26__leaf_clk),
    .X(clknet_leaf_81_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1647 (.A(_02692_),
    .X(net1647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1648 (.A(_02345_),
    .X(net1648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1669 (.A(_01844_),
    .X(net1669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_89_clk (.A(clknet_5_24__leaf_clk),
    .X(clknet_leaf_89_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1650 (.A(_01935_),
    .X(net1650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1655 (.A(_05136_),
    .X(net1655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1660 (.A(_01905_),
    .X(net1660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_63_clk (.A(clknet_5_29__leaf_clk),
    .X(clknet_leaf_63_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_55_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_55_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_73_clk (.A(clknet_5_31__leaf_clk),
    .X(clknet_leaf_73_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1659 (.A(_02338_),
    .X(net1659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1662 (.A(_04105_),
    .X(net1662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_58_clk (.A(clknet_5_30__leaf_clk),
    .X(clknet_leaf_58_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_53_clk (.A(clknet_5_18__leaf_clk),
    .X(clknet_leaf_53_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1678 (.A(net1677),
    .X(net1678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1676 (.A(_06962_),
    .X(net1676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_48_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1686 (.A(_01840_),
    .X(net1686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_45_clk (.A(clknet_5_22__leaf_clk),
    .X(clknet_leaf_45_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_5_20__leaf_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_5_23__leaf_clk),
    .X(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1690 (.A(_03828_),
    .X(net1690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1673 (.A(_04460_),
    .X(net1673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1819 (.A(\acc_sum.reg2en.q[0] ),
    .X(net1819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_5_19__leaf_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1685 (.A(_01871_),
    .X(net1685),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1677 (.A(_06962_),
    .X(net1677),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_5_17__leaf_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1688 (.A(_04076_),
    .X(net1688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_5_16__leaf_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1687 (.A(_01840_),
    .X(net1687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_5_5__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1721 (.A(_07076_),
    .X(net1721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1700 (.A(_06837_),
    .X(net1700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout140 (.A(net141),
    .X(net140),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout139 (.A(net140),
    .X(net139),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout138 (.A(net139),
    .X(net138),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout131 (.A(net140),
    .X(net131),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1714 (.A(net1713),
    .X(net1714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1718 (.A(_02650_),
    .X(net1718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1705 (.A(_02654_),
    .X(net1705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1706 (.A(_02654_),
    .X(net1706),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1693 (.A(_07055_),
    .X(net1693),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout128 (.A(net141),
    .X(net128),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout122 (.A(net128),
    .X(net122),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1710 (.A(_04654_),
    .X(net1710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1711 (.A(_02578_),
    .X(net1711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1712 (.A(_06907_),
    .X(net1712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1730 (.A(_06571_),
    .X(net1730),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout112 (.A(net113),
    .X(net112),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout111 (.A(net113),
    .X(net111),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1727 (.A(_05583_),
    .X(net1727),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1717 (.A(_06574_),
    .X(net1717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1723 (.A(_07027_),
    .X(net1723),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1726 (.A(net1725),
    .X(net1726),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1732 (.A(_06559_),
    .X(net1732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1733 (.A(net1732),
    .X(net1733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1757 (.A(_05498_),
    .X(net1757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout102 (.A(net104),
    .X(net102),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout101 (.A(net102),
    .X(net101),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1734 (.A(_06366_),
    .X(net1734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout98 (.A(net100),
    .X(net98),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1762 (.A(net1761),
    .X(net1762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1740 (.A(_02726_),
    .X(net1740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1742 (.A(_02569_),
    .X(net1742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout87 (.A(net88),
    .X(net87),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1747 (.A(_02058_),
    .X(net1747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1748 (.A(_01756_),
    .X(net1748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout83 (.A(net86),
    .X(net83),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout80 (.A(net81),
    .X(net80),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1746 (.A(_04073_),
    .X(net1746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1768 (.A(_03782_),
    .X(net1768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1780 (.A(net1779),
    .X(net1780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout73 (.A(net74),
    .X(net73),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1894 (.A(net1893),
    .X(net1894),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1817 (.A(net1816),
    .X(net1817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1766 (.A(_03988_),
    .X(net1766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1758 (.A(net1757),
    .X(net1758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout66 (.A(net67),
    .X(net66),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1782 (.A(_01779_),
    .X(net1782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1794 (.A(\acc_sub.exp_mant_logic0.b[6] ),
    .X(net1794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1765 (.A(_03988_),
    .X(net1765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1795 (.A(\acc_sub.exp_mant_logic0.b[5] ),
    .X(net1795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1804 (.A(net1802),
    .X(net1804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1771 (.A(_03359_),
    .X(net1771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1784 (.A(net1783),
    .X(net1784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1785 (.A(_01490_),
    .X(net1785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1798 (.A(net1797),
    .X(net1798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1770 (.A(_03361_),
    .X(net1770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout54 (.A(net55),
    .X(net54),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout53 (.A(net55),
    .X(net53),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1773 (.A(_02965_),
    .X(net1773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1791 (.A(net1790),
    .X(net1791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1781 (.A(net1779),
    .X(net1781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1783 (.A(_01492_),
    .X(net1783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1787 (.A(\acc_sub.seg_reg1.q[21] ),
    .X(net1787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1807 (.A(\acc_sum.add_renorm0.mantisa[11] ),
    .X(net1807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1789 (.A(net1788),
    .X(net1789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout47 (.A(net72),
    .X(net47),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1803 (.A(net1802),
    .X(net1803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1850 (.A(\fp16_sum_pipe.reg3en.q[0] ),
    .X(net1850),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1778 (.A(net1777),
    .X(net1778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1800 (.A(\acc_sub.reg3en.q[0] ),
    .X(net1800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1806 (.A(net1805),
    .X(net1806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1827 (.A(\fp16_res_pipe.exp_mant_logic0.a[6] ),
    .X(net1827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1805 (.A(\acc_sum.add_renorm0.mantisa[11] ),
    .X(net1805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1796 (.A(\acc_sub.reg1en.q[0] ),
    .X(net1796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout41 (.A(net42),
    .X(net41),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout43 (.A(net46),
    .X(net43),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout42 (.A(net47),
    .X(net42),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout44 (.A(net46),
    .X(net44),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1797 (.A(\acc_sub.reg2en.q[0] ),
    .X(net1797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout40 (.A(net41),
    .X(net40),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1801 (.A(\acc_sub.reg3en.q[0] ),
    .X(net1801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1802 (.A(\acc_sum.seg_reg1.q[21] ),
    .X(net1802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1907 (.A(load_en),
    .X(net1907),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1849 (.A(net1848),
    .X(net1849),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1815 (.A(net1814),
    .X(net1815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1808 (.A(\acc_sum.exp_mant_logic0.a[6] ),
    .X(net1808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1848 (.A(net1847),
    .X(net1848),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1809 (.A(\acc_sum.exp_mant_logic0.a[5] ),
    .X(net1809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1862 (.A(\fpmul.reg2en.q[0] ),
    .X(net1862),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1810 (.A(\acc_sum.exp_mant_logic0.a[4] ),
    .X(net1810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1823 (.A(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .X(net1823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1847 (.A(\fp16_sum_pipe.reg2en.q[0] ),
    .X(net1847),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1840 (.A(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .X(net1840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1841 (.A(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .X(net1841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1811 (.A(\acc_sum.exp_mant_logic0.b[6] ),
    .X(net1811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1833 (.A(net1832),
    .X(net1833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1846 (.A(net1845),
    .X(net1846),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1812 (.A(\acc_sum.exp_mant_logic0.b[5] ),
    .X(net1812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1875 (.A(\fpmul.reg1en.q[0] ),
    .X(net1875),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1813 (.A(\acc_sum.reg1en.q[0] ),
    .X(net1813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1814 (.A(\acc_sum.reg2en.q[0] ),
    .X(net1814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1826 (.A(\fp16_res_pipe.add_renorm0.mantisa[11] ),
    .X(net1826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1834 (.A(net1833),
    .X(net1834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1828 (.A(\fp16_res_pipe.exp_mant_logic0.a[5] ),
    .X(net1828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1829 (.A(\fp16_res_pipe.exp_mant_logic0.b[6] ),
    .X(net1829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1835 (.A(\fp16_res_pipe.reg3en.q[0] ),
    .X(net1835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1853 (.A(\fpmul.seg_reg0.q[15] ),
    .X(net1853),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1830 (.A(\fp16_res_pipe.exp_mant_logic0.b[5] ),
    .X(net1830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout38 (.A(net39),
    .X(net38),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout36 (.A(net38),
    .X(net36),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout37 (.A(net38),
    .X(net37),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout39 (.A(net72),
    .X(net39),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1836 (.A(\fp16_sum_pipe.seg_reg1.q[21] ),
    .X(net1836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1873 (.A(\fpmul.reg1en.q[0] ),
    .X(net1873),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1901 (.A(net1900),
    .X(net1901),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1845 (.A(net1844),
    .X(net1845),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1839 (.A(net1838),
    .X(net1839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1831 (.A(\fp16_res_pipe.reg1en.q[0] ),
    .X(net1831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1893 (.A(\acc_sub.reg1en.d[0] ),
    .X(net1893),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout34 (.A(net39),
    .X(net34),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1852 (.A(net1851),
    .X(net1852),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout33 (.A(net34),
    .X(net33),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout35 (.A(net38),
    .X(net35),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1832 (.A(\fp16_res_pipe.reg2en.q[0] ),
    .X(net1832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1837 (.A(net1836),
    .X(net1837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1838 (.A(\fp16_sum_pipe.add_renorm0.mantisa[11] ),
    .X(net1838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1872 (.A(net1871),
    .X(net1872),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1842 (.A(\fp16_sum_pipe.exp_mant_logic0.b[5] ),
    .X(net1842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1871 (.A(net1870),
    .X(net1871),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1843 (.A(\fp16_sum_pipe.reg1en.q[0] ),
    .X(net1843),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1854 (.A(\fpmul.reg_a_out[6] ),
    .X(net1854),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1917 (.A(net1916),
    .X(net1917),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1892 (.A(net1891),
    .X(net1892),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1844 (.A(\fp16_sum_pipe.reg2en.q[0] ),
    .X(net1844),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1874 (.A(net1873),
    .X(net1874),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1905 (.A(net1903),
    .X(net1905),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1900 (.A(net1897),
    .X(net1900),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1890 (.A(net1889),
    .X(net1890),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1915 (.A(net1913),
    .X(net1915),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1855 (.A(\fpmul.reg_a_out[5] ),
    .X(net1855),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1913 (.A(net1912),
    .X(net1913),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1912 (.A(net1911),
    .X(net1912),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1902 (.A(net1900),
    .X(net1902),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1914 (.A(net1913),
    .X(net1914),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1891 (.A(net1889),
    .X(net1891),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1923 (.A(net1922),
    .X(net1923),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1932 (.A(net1930),
    .X(net1932),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout6 (.A(net15),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(rst),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1909 (.A(\fp16_res_pipe.reg1en.d[0] ),
    .X(net1909),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1945 (.A(net1944),
    .X(net1945),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1910 (.A(\fp16_res_pipe.reg1en.d[0] ),
    .X(net1910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1953 (.A(net1952),
    .X(net1953),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1856 (.A(\fpmul.reg_a_out[4] ),
    .X(net1856),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1899 (.A(net1898),
    .X(net1899),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1857 (.A(\fpmul.reg_a_out[3] ),
    .X(net1857),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1858 (.A(\fpmul.reg_a_out[2] ),
    .X(net1858),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout16 (.A(net17),
    .X(net16),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1931 (.A(net1930),
    .X(net1931),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1859 (.A(\fpmul.reg_a_out[1] ),
    .X(net1859),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1860 (.A(\fpmul.reg_a_out[0] ),
    .X(net1860),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1861 (.A(\fpmul.reg2en.q[0] ),
    .X(net1861),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1863 (.A(\fpmul.reg_b_out[6] ),
    .X(net1863),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1864 (.A(\fpmul.reg_b_out[5] ),
    .X(net1864),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1866 (.A(\fpmul.reg_b_out[3] ),
    .X(net1866),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1865 (.A(\fpmul.reg_b_out[4] ),
    .X(net1865),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1950 (.A(net1948),
    .X(net1950),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout17 (.A(net18),
    .X(net17),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1867 (.A(\fpmul.reg_b_out[2] ),
    .X(net1867),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1928 (.A(net1927),
    .X(net1928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1868 (.A(\fpmul.reg_b_out[1] ),
    .X(net1868),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1930 (.A(net1924),
    .X(net1930),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1869 (.A(\fpmul.reg_b_out[0] ),
    .X(net1869),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1929 (.A(net1928),
    .X(net1929),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1870 (.A(\fpmul.reg1en.q[0] ),
    .X(net1870),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1920 (.A(net1912),
    .X(net1920),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1925 (.A(net1924),
    .X(net1925),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1946 (.A(net1944),
    .X(net1946),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1927 (.A(net1925),
    .X(net1927),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1952 (.A(net1951),
    .X(net1952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1933 (.A(net1930),
    .X(net1933),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1937 (.A(\fpdiv.reg1en.d[0] ),
    .X(net1937),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1942 (.A(net1941),
    .X(net1942),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1938 (.A(\fpdiv.reg1en.d[0] ),
    .X(net1938),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1939 (.A(net1938),
    .X(net1939),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1934 (.A(net1933),
    .X(net1934),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1940 (.A(net1939),
    .X(net1940),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout31 (.A(net39),
    .X(net31),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1944 (.A(\fpdiv.reg1en.d[0] ),
    .X(net1944),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1941 (.A(\fpdiv.reg1en.d[0] ),
    .X(net1941),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout30 (.A(net31),
    .X(net30),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout26 (.A(net28),
    .X(net26),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout27 (.A(net28),
    .X(net27),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout29 (.A(net30),
    .X(net29),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout28 (.A(net31),
    .X(net28),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout32 (.A(net34),
    .X(net32),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1943 (.A(net1941),
    .X(net1943),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1951 (.A(\fpmul.reg1en.d[0] ),
    .X(net1951),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1959 (.A(net1958),
    .X(net1959),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1956 (.A(net1954),
    .X(net1956),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1949 (.A(net1948),
    .X(net1949),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout15 (.A(net72),
    .X(net15),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1958 (.A(\fpmul.reg1en.d[0] ),
    .X(net1958),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1962 (.A(net1961),
    .X(net1962),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1954 (.A(\fpmul.reg1en.d[0] ),
    .X(net1954),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1961 (.A(\fpmul.reg1en.d[0] ),
    .X(net1961),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout25 (.A(net28),
    .X(net25),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout7 (.A(net15),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout10 (.A(net15),
    .X(net10),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1957 (.A(net1954),
    .X(net1957),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1960 (.A(net1959),
    .X(net1960),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout9 (.A(net10),
    .X(net9),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input1 (.A(mosi),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 input3 (.A(ss),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout11 (.A(net13),
    .X(net11),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1667 (.A(net1666),
    .X(net1667),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout8 (.A(net15),
    .X(net8),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout14 (.A(net15),
    .X(net14),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout13 (.A(net14),
    .X(net13),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout12 (.A(net13),
    .X(net12),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output4 (.A(net4),
    .X(miso),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1679 (.A(_06962_),
    .X(net1679),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1955 (.A(net1954),
    .X(net1955),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1656 (.A(net1655),
    .X(net1656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1666 (.A(net1665),
    .X(net1666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1921 (.A(net1920),
    .X(net1921),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1879 (.A(net1877),
    .X(net1879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1634 (.A(_05256_),
    .X(net1634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1882 (.A(net1881),
    .X(net1882),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1884 (.A(net1883),
    .X(net1884),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout23 (.A(net24),
    .X(net23),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1883 (.A(net1882),
    .X(net1883),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1878 (.A(net1877),
    .X(net1878),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1880 (.A(\fpmul.reg1en.q[0] ),
    .X(net1880),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1877 (.A(net1875),
    .X(net1877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1881 (.A(net1880),
    .X(net1881),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout24 (.A(net39),
    .X(net24),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1702 (.A(net1701),
    .X(net1702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1922 (.A(\fp16_sum_pipe.reg1en.d[0] ),
    .X(net1922),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1697 (.A(_05075_),
    .X(net1697),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1668 (.A(_02865_),
    .X(net1668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1825 (.A(net1824),
    .X(net1825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1822 (.A(\fp16_res_pipe.seg_reg1.q[21] ),
    .X(net1822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout21 (.A(net23),
    .X(net21),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1779 (.A(_01779_),
    .X(net1779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout20 (.A(net24),
    .X(net20),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1675 (.A(_03453_),
    .X(net1675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1799 (.A(net1797),
    .X(net1799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1635 (.A(_05151_),
    .X(net1635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout19 (.A(net24),
    .X(net19),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1786 (.A(net1785),
    .X(net1786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1680 (.A(_05052_),
    .X(net1680),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1696 (.A(_07055_),
    .X(net1696),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout18 (.A(net24),
    .X(net18),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout22 (.A(net23),
    .X(net22),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1897 (.A(\acc_sum.reg1en.d[0] ),
    .X(net1897),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1935 (.A(net1923),
    .X(net1935),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1729 (.A(net1728),
    .X(net1729),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1720 (.A(_07076_),
    .X(net1720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1695 (.A(net1693),
    .X(net1695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1681 (.A(_05049_),
    .X(net1681),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1636 (.A(_04272_),
    .X(net1636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1948 (.A(net1944),
    .X(net1948),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1896 (.A(\acc_sum.reg1en.d[0] ),
    .X(net1896),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1777 (.A(net1774),
    .X(net1777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1924 (.A(net1923),
    .X(net1924),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1898 (.A(net1897),
    .X(net1898),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1926 (.A(net1925),
    .X(net1926),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1947 (.A(net1946),
    .X(net1947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1903 (.A(net1902),
    .X(net1903),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1904 (.A(net1903),
    .X(net1904),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1936 (.A(net1935),
    .X(net1936),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1699 (.A(_03146_),
    .X(net1699),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1637 (.A(_04150_),
    .X(net1637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1682 (.A(_04056_),
    .X(net1682),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1895 (.A(net1893),
    .X(net1895),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1911 (.A(net1910),
    .X(net1911),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1908 (.A(load_en),
    .X(net1908),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1906 (.A(net1902),
    .X(net1906),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout5 (.A(net6),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1820 (.A(\acc_sum.reg3en.q[0] ),
    .X(net1820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1889 (.A(net1885),
    .X(net1889),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1887 (.A(net1886),
    .X(net1887),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1888 (.A(net1887),
    .X(net1888),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 place1886 (.A(net1885),
    .X(net1886),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1885 (.A(\acc_sub.reg1en.d[0] ),
    .X(net1885),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1919 (.A(net1912),
    .X(net1919),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 place1638 (.A(_02475_),
    .X(net1638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_103_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_103_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_104_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_104_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_105_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_105_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_106_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_106_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_107_clk (.A(clknet_5_14__leaf_clk),
    .X(clknet_leaf_107_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_108_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_108_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_109_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_109_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_110_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_110_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_111_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_111_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_112_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_112_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_114_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_114_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_115_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_115_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_116_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_116_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_117_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_117_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_118_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_118_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_119_clk (.A(clknet_5_10__leaf_clk),
    .X(clknet_leaf_119_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_120_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_120_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_121_clk (.A(clknet_5_11__leaf_clk),
    .X(clknet_leaf_121_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_122_clk (.A(clknet_5_9__leaf_clk),
    .X(clknet_leaf_122_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_123_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_123_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_124_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_124_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_125_clk (.A(clknet_5_12__leaf_clk),
    .X(clknet_leaf_125_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_126_clk (.A(clknet_5_13__leaf_clk),
    .X(clknet_leaf_126_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_127_clk (.A(clknet_5_7__leaf_clk),
    .X(clknet_leaf_127_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_128_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_128_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_129_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_129_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_130_clk (.A(clknet_5_6__leaf_clk),
    .X(clknet_leaf_130_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_131_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_131_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_132_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_132_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_134_clk (.A(clknet_5_3__leaf_clk),
    .X(clknet_leaf_134_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_135_clk (.A(clknet_5_8__leaf_clk),
    .X(clknet_leaf_135_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_136_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_136_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_137_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_137_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_139_clk (.A(clknet_5_2__leaf_clk),
    .X(clknet_leaf_139_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_140_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_140_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_141_clk (.A(clknet_5_1__leaf_clk),
    .X(clknet_leaf_141_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_142_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_142_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_143_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_143_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_144_clk (.A(clknet_5_0__leaf_clk),
    .X(clknet_leaf_144_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_0_0_clk (.A(clknet_0_clk),
    .X(clknet_4_0_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_1_0_clk (.A(clknet_0_clk),
    .X(clknet_4_1_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_2_0_clk (.A(clknet_0_clk),
    .X(clknet_4_2_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_3_0_clk (.A(clknet_0_clk),
    .X(clknet_4_3_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_4_0_clk (.A(clknet_0_clk),
    .X(clknet_4_4_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_5_0_clk (.A(clknet_0_clk),
    .X(clknet_4_5_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_6_0_clk (.A(clknet_0_clk),
    .X(clknet_4_6_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_7_0_clk (.A(clknet_0_clk),
    .X(clknet_4_7_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_8_0_clk (.A(clknet_0_clk),
    .X(clknet_4_8_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_9_0_clk (.A(clknet_0_clk),
    .X(clknet_4_9_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_10_0_clk (.A(clknet_0_clk),
    .X(clknet_4_10_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_11_0_clk (.A(clknet_0_clk),
    .X(clknet_4_11_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_12_0_clk (.A(clknet_0_clk),
    .X(clknet_4_12_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_13_0_clk (.A(clknet_0_clk),
    .X(clknet_4_13_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_14_0_clk (.A(clknet_0_clk),
    .X(clknet_4_14_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_4_15_0_clk (.A(clknet_0_clk),
    .X(clknet_4_15_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_0__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_1__f_clk (.A(clknet_4_0_0_clk),
    .X(clknet_5_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_2__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_3__f_clk (.A(clknet_4_1_0_clk),
    .X(clknet_5_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_4__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_5__f_clk (.A(clknet_4_2_0_clk),
    .X(clknet_5_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_6__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_7__f_clk (.A(clknet_4_3_0_clk),
    .X(clknet_5_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_8__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_8__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_9__f_clk (.A(clknet_4_4_0_clk),
    .X(clknet_5_9__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_10__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_10__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_11__f_clk (.A(clknet_4_5_0_clk),
    .X(clknet_5_11__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_12__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_12__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_13__f_clk (.A(clknet_4_6_0_clk),
    .X(clknet_5_13__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_14__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_14__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_15__f_clk (.A(clknet_4_7_0_clk),
    .X(clknet_5_15__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_16__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_16__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_17__f_clk (.A(clknet_4_8_0_clk),
    .X(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_18__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_18__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_19__f_clk (.A(clknet_4_9_0_clk),
    .X(clknet_5_19__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_20__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_20__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_21__f_clk (.A(clknet_4_10_0_clk),
    .X(clknet_5_21__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_22__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_22__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_23__f_clk (.A(clknet_4_11_0_clk),
    .X(clknet_5_23__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_24__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_24__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_25__f_clk (.A(clknet_4_12_0_clk),
    .X(clknet_5_25__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_26__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_26__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_27__f_clk (.A(clknet_4_13_0_clk),
    .X(clknet_5_27__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_28__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_28__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_29__f_clk (.A(clknet_4_14_0_clk),
    .X(clknet_5_29__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_30__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_30__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_5_31__f_clk (.A(clknet_4_15_0_clk),
    .X(clknet_5_31__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload0 (.A(clknet_5_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload1 (.VDD(VPWR),
    .A(clknet_5_3__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_5_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload3 (.A(clknet_5_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload4 (.VDD(VPWR),
    .A(clknet_5_9__leaf_clk),
    .VSS(VGND));
 sg13g2_buf_8 clkload5 (.A(clknet_5_11__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload6 (.A(clknet_5_13__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload7 (.A(clknet_5_15__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload8 (.A(clknet_5_17__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload9 (.A(clknet_5_19__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload10 (.A(clknet_5_21__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload11 (.A(clknet_5_23__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload12 (.A(clknet_5_25__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload13 (.A(clknet_5_27__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload14 (.A(clknet_5_29__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload15 (.A(clknet_5_31__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload16 (.A(clknet_leaf_140_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload17 (.A(clknet_leaf_143_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload18 (.A(clknet_leaf_144_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload19 (.A(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload20 (.A(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload21 (.VDD(VPWR),
    .A(clknet_leaf_2_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload22 (.A(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload23 (.A(clknet_leaf_136_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload24 (.VDD(VPWR),
    .A(clknet_leaf_137_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload25 (.VDD(VPWR),
    .A(clknet_leaf_139_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload26 (.VDD(VPWR),
    .A(clknet_leaf_129_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload27 (.VDD(VPWR),
    .A(clknet_leaf_131_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload28 (.A(clknet_leaf_134_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload29 (.A(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload30 (.VDD(VPWR),
    .A(clknet_leaf_8_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload31 (.A(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload32 (.A(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload33 (.A(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload34 (.A(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload35 (.A(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload36 (.VDD(VPWR),
    .A(clknet_leaf_12_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload37 (.A(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload38 (.VDD(VPWR),
    .A(clknet_leaf_16_clk),
    .VSS(VGND));
 sg13g2_inv_1 clkload39 (.VDD(VPWR),
    .A(clknet_leaf_15_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload40 (.A(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload41 (.A(clknet_leaf_114_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload42 (.A(clknet_leaf_116_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload43 (.A(clknet_leaf_135_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload44 (.A(clknet_leaf_117_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload45 (.A(clknet_leaf_118_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload46 (.A(clknet_leaf_122_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload47 (.A(clknet_leaf_108_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload48 (.A(clknet_leaf_109_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload49 (.A(clknet_leaf_110_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload50 (.A(clknet_leaf_111_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload51 (.A(clknet_leaf_98_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload52 (.A(clknet_leaf_120_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload53 (.A(clknet_leaf_92_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload54 (.A(clknet_leaf_93_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload55 (.A(clknet_leaf_96_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload56 (.A(clknet_leaf_124_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload57 (.A(clknet_leaf_94_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload58 (.A(clknet_leaf_95_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload59 (.A(clknet_leaf_126_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload60 (.A(clknet_leaf_103_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 clkload61 (.A(clknet_leaf_105_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload62 (.A(clknet_leaf_106_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload63 (.VDD(VPWR),
    .A(clknet_leaf_107_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload64 (.A(clknet_leaf_100_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload65 (.A(clknet_leaf_101_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload66 (.A(clknet_leaf_102_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload67 (.A(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload68 (.A(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload69 (.A(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload70 (.VDD(VPWR),
    .A(clknet_leaf_30_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload71 (.A(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload72 (.A(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload73 (.A(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload74 (.A(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload75 (.VDD(VPWR),
    .A(clknet_leaf_21_clk),
    .VSS(VGND));
 sg13g2_inv_2 clkload76 (.A(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload77 (.A(clknet_leaf_52_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload78 (.A(clknet_leaf_55_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload79 (.A(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload80 (.A(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload81 (.A(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload82 (.A(clknet_leaf_48_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload83 (.A(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload84 (.A(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload85 (.A(clknet_leaf_47_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload86 (.VDD(VPWR),
    .A(clknet_leaf_49_clk),
    .VSS(VGND));
 sg13g2_inv_8 clkload87 (.A(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload88 (.VDD(VPWR),
    .A(clknet_leaf_42_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload89 (.A(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload90 (.A(clknet_leaf_82_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload91 (.A(clknet_leaf_88_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload92 (.A(clknet_leaf_89_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload93 (.A(clknet_leaf_90_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload94 (.A(clknet_leaf_57_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload95 (.A(clknet_leaf_85_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload96 (.VDD(VPWR),
    .A(clknet_leaf_86_clk),
    .VSS(VGND));
 sg13g2_buf_1 clkload97 (.A(clknet_leaf_78_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload98 (.A(clknet_leaf_79_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload99 (.VDD(VPWR),
    .A(clknet_leaf_80_clk),
    .VSS(VGND));
 sg13g2_inv_4 clkload100 (.A(clknet_leaf_83_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload101 (.A(clknet_leaf_75_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload102 (.A(clknet_leaf_76_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload103 (.A(clknet_leaf_77_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload104 (.A(clknet_leaf_61_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload105 (.A(clknet_leaf_62_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload106 (.A(clknet_leaf_68_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload107 (.A(clknet_leaf_66_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload108 (.A(clknet_leaf_59_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload109 (.A(clknet_leaf_70_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload110 (.A(clknet_leaf_72_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload111 (.A(clknet_leaf_74_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload112 (.VDD(VPWR),
    .A(clknet_leaf_67_clk),
    .VSS(VGND));
 sg13g2_inv_8 clkload113 (.A(clknet_leaf_71_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 clkload114 (.A(clknet_leaf_73_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_50_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_50_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_50_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_50_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_51_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_51_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_51_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_51_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_52_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_52_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_52_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_52_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_53_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_53_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_53_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_53_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_54_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_54_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_54_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_54_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_55_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_55_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_55_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_55_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_56_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_56_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_56_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_56_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_57_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_57_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_57_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_57_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_58_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_58_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_58_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_58_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_59_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_59_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_59_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_59_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_60_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_60_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_60_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_60_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_61_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_61_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_61_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_61_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_62_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_62_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_62_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_62_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_63_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_63_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_63_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_63_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_64_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_64_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_64_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_64_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_65_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_65_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_65_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_65_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_66_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_66_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_66_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_66_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_67_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_67_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_67_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_67_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_68_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_68_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_68_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_68_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_69_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_69_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_69_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_69_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_70_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_70_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_70_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_70_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_71_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_71_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_71_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_71_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_34 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_41 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_72_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_72_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_72_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_72_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_73_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_73_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_73_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_73_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_74_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_74_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_74_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_74_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_227 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_75_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_75_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_75_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_75_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_76_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_76_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_76_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_76_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_77_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_77_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_77_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_77_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_78_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_78_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_78_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_78_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_79_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_79_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_79_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_79_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_80_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_80_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_80_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_80_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_6 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_81_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_81_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_81_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_81_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_82_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_82_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_82_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_82_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_83_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_83_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_83_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_83_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_84_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_84_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_84_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_84_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_85_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_85_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_85_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_85_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_86_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_86_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_86_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_86_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_87_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_87_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_87_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_87_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_88_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_88_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_88_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_88_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_170 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_89_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_89_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_89_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_89_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_90_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_90_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_90_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_90_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_177 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_91_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_91_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_91_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_91_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_92_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_92_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_92_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_92_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_93_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_93_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_93_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_93_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_94_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_94_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_94_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_94_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_95_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_95_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_95_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_95_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_96_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_96_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_96_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_96_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_97_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_97_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_97_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_97_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_98_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_98_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_98_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_98_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_99_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_99_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_99_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_99_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_100_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_100_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_100_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_100_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_101_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_101_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_101_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_101_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_102_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_102_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_102_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_102_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_108 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_589 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_103_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_103_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_103_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_103_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_31 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_104_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_104_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_104_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_104_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_105_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_105_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_105_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_105_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_23 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_158 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_172 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_389 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_106_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_106_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_106_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_106_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_279 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_107_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_107_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_107_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_107_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_108_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_108_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_108_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_108_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_144 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_109_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_109_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_109_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_109_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_110_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_110_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_110_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_110_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_288 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_111_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_111_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_111_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_111_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_169 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_112_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_112_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_112_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_112_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_596 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_112_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_112_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_112_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_112_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_113_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_113_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_113_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_113_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_114_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_114_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_114_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_114_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_114_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_114_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_114_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_114_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_114_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_115_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_115_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_115_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_115_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_115_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_610 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_115_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_115_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_115_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_115_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_5 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_12 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_33 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_54 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_131 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_116_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_116_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_116_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_116_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_116_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_116_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_116_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_117_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_368 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_117_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_117_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_117_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_117_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_117_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_117_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_424 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_118_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_118_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_118_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_118_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_119_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_277 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_119_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_119_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_119_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_119_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_119_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_119_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_119_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_119_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_503 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_120_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_120_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_120_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_120_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_121_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_121_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_121_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_121_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_122_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_122_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_122_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_122_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_123_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_123_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_123_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_123_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_124_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_124_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_124_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_124_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_124_653 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_124_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_124_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_124_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_125_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_125_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_125_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_125_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_125_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_125_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_125_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_125_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_126_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_126_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_126_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_126_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_49 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_287 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_308 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_329 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_127_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_127_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_458 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_127_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_127_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_478 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_485 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_127_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_679 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_127_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_127_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_127_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_127_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_127_1013 (.VDD(VPWR),
    .VSS(VGND));
endmodule
