* NGSPICE file created from bfloat16_spi_top.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nor4_2 abstract view
.subckt sg13g2_nor4_2 A B C Y VSS VDD D
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

.subckt bfloat16_spi_top VGND VPWR clk miso mosi rst ss
XFILLER_79_380 VPWR VGND sg13g2_fill_2
XFILLER_95_873 VPWR VGND sg13g2_fill_1
X_09671_ _03787_ VPWR _01240_ VGND _02729_ _03785_ sg13g2_o21ai_1
XFILLER_55_726 VPWR VGND sg13g2_fill_1
XFILLER_55_704 VPWR VGND sg13g2_decap_8
XFILLER_54_203 VPWR VGND sg13g2_decap_8
XFILLER_94_383 VPWR VGND sg13g2_fill_1
X_08622_ _02792_ _02759_ _02782_ _02745_ _02844_ VPWR VGND sg13g2_and4_1
X_08553_ acc_sum.op_sign_logic0.mantisa_b\[5\] _02776_ _02777_ VPWR VGND sg13g2_nor2_1
XFILLER_82_578 VPWR VGND sg13g2_fill_1
XFILLER_82_556 VPWR VGND sg13g2_decap_8
XFILLER_54_269 VPWR VGND sg13g2_fill_1
XFILLER_36_962 VPWR VGND sg13g2_decap_8
X_07504_ _01826_ _01825_ acc_sub.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
X_08484_ _02712_ VPWR _02713_ VGND fpdiv.divider0.remainder_reg\[6\] _02692_ sg13g2_o21ai_1
XFILLER_70_729 VPWR VGND sg13g2_decap_8
XFILLER_35_483 VPWR VGND sg13g2_decap_8
XFILLER_23_601 VPWR VGND sg13g2_decap_8
X_07435_ fpdiv.divider0.divisor_reg\[8\] net1750 _01767_ VPWR VGND sg13g2_nor2_1
XFILLER_35_1009 VPWR VGND sg13g2_decap_4
XFILLER_23_634 VPWR VGND sg13g2_fill_2
XFILLER_51_976 VPWR VGND sg13g2_fill_2
XFILLER_22_155 VPWR VGND sg13g2_fill_2
X_07366_ _01720_ net1799 acc_sub.seg_reg0.q\[24\] VPWR VGND sg13g2_nand2_1
XFILLER_10_328 VPWR VGND sg13g2_fill_2
X_07297_ _01663_ VPWR _01483_ VGND _01656_ _01661_ sg13g2_o21ai_1
X_09105_ _03100_ VPWR _03287_ VGND _03194_ _03286_ sg13g2_o21ai_1
XFILLER_108_216 VPWR VGND sg13g2_fill_1
X_09036_ net1790 _03170_ _03221_ _03222_ VPWR VGND sg13g2_a21o_1
XFILLER_116_271 VPWR VGND sg13g2_decap_8
XFILLER_105_923 VPWR VGND sg13g2_decap_8
XFILLER_89_100 VPWR VGND sg13g2_fill_2
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_120_904 VPWR VGND sg13g2_decap_8
XFILLER_117_77 VPWR VGND sg13g2_decap_8
XFILLER_77_26 VPWR VGND sg13g2_decap_8
XFILLER_2_549 VPWR VGND sg13g2_fill_2
XFILLER_89_166 VPWR VGND sg13g2_decap_4
XFILLER_77_317 VPWR VGND sg13g2_decap_8
X_09938_ VPWR _04034_ fp16_res_pipe.exp_mant_logic0.b\[8\] VGND sg13g2_inv_1
X_09869_ _03975_ _03687_ _03655_ VPWR VGND sg13g2_nand2_1
XFILLER_19_929 VPWR VGND sg13g2_decap_8
X_12880_ _06658_ _06657_ net1732 VPWR VGND sg13g2_nand2_1
X_11900_ _05780_ VPWR _01004_ VGND net1877 _05779_ sg13g2_o21ai_1
XFILLER_46_748 VPWR VGND sg13g2_fill_2
XFILLER_45_225 VPWR VGND sg13g2_decap_8
X_11831_ _01023_ _05729_ _05730_ VPWR VGND sg13g2_nand2_1
XFILLER_45_258 VPWR VGND sg13g2_decap_8
X_14550_ _00351_ VGND VPWR _01086_ acc_sum.op_sign_logic0.mantisa_a\[2\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
XFILLER_54_792 VPWR VGND sg13g2_fill_1
XFILLER_26_63 VPWR VGND sg13g2_decap_8
XFILLER_27_995 VPWR VGND sg13g2_decap_8
X_13501_ VPWR _00052_ net84 VGND sg13g2_inv_1
XFILLER_13_111 VPWR VGND sg13g2_decap_8
X_11762_ fp16_sum_pipe.add_renorm0.exp\[1\] _05665_ _05536_ _05666_ VPWR VGND sg13g2_nand3_1
X_14481_ _00282_ VGND VPWR _01019_ add_result\[6\] clknet_leaf_100_clk sg13g2_dfrbpq_1
XFILLER_13_155 VPWR VGND sg13g2_decap_8
X_10713_ VPWR _04726_ _04724_ VGND sg13g2_inv_1
X_13432_ _07095_ net1720 instr\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_9_126 VPWR VGND sg13g2_decap_8
X_10644_ _04657_ _04650_ _04656_ VPWR VGND sg13g2_nand2_1
XFILLER_42_84 VPWR VGND sg13g2_decap_8
X_10575_ _04600_ VPWR _01149_ VGND net1926 _02197_ sg13g2_o21ai_1
XFILLER_6_800 VPWR VGND sg13g2_fill_1
X_12314_ _06160_ net1857 net1867 VPWR VGND sg13g2_nand2_2
XFILLER_10_884 VPWR VGND sg13g2_decap_8
XFILLER_127_569 VPWR VGND sg13g2_decap_8
X_13294_ VPWR VGND acc_sub.y\[4\] _07007_ net1711 net1728 _07008_ acc_sum.y\[4\] sg13g2_a221oi_1
X_12245_ _06072_ _06074_ _06091_ VPWR VGND sg13g2_nor2_1
XFILLER_6_899 VPWR VGND sg13g2_decap_8
XFILLER_123_764 VPWR VGND sg13g2_decap_8
XFILLER_96_604 VPWR VGND sg13g2_decap_8
X_12176_ VPWR _06022_ _06005_ VGND sg13g2_inv_1
XFILLER_122_252 VPWR VGND sg13g2_decap_8
XFILLER_111_915 VPWR VGND sg13g2_decap_8
XFILLER_110_403 VPWR VGND sg13g2_decap_8
XFILLER_69_829 VPWR VGND sg13g2_decap_8
X_11127_ VGND VPWR _05046_ _05082_ _05097_ _05096_ sg13g2_a21oi_1
XFILLER_3_56 VPWR VGND sg13g2_decap_8
XFILLER_95_147 VPWR VGND sg13g2_decap_8
XFILLER_77_862 VPWR VGND sg13g2_fill_1
X_11058_ _04998_ _05010_ _05036_ VPWR VGND sg13g2_nor2_1
X_10009_ _04097_ _04096_ _03993_ VPWR VGND sg13g2_nand2_1
X_14817_ _00618_ VGND VPWR _01341_ acc_sum.add_renorm0.mantisa\[6\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_36_247 VPWR VGND sg13g2_decap_8
XFILLER_18_962 VPWR VGND sg13g2_decap_8
XFILLER_91_375 VPWR VGND sg13g2_decap_4
XFILLER_51_217 VPWR VGND sg13g2_fill_1
XFILLER_33_932 VPWR VGND sg13g2_decap_8
XFILLER_17_472 VPWR VGND sg13g2_decap_8
X_14748_ _00549_ VGND VPWR _01276_ fp16_res_pipe.add_renorm0.mantisa\[11\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_2
XFILLER_32_420 VPWR VGND sg13g2_decap_8
XFILLER_20_615 VPWR VGND sg13g2_fill_1
X_14679_ _00480_ VGND VPWR _01207_ fp16_res_pipe.op_sign_logic0.mantisa_a\[5\] clknet_leaf_144_clk
+ sg13g2_dfrbpq_2
XFILLER_20_637 VPWR VGND sg13g2_decap_4
XFILLER_121_1012 VPWR VGND sg13g2_fill_2
XFILLER_121_1001 VPWR VGND sg13g2_decap_8
X_07151_ VPWR _01523_ acc_sub.op_sign_logic0.mantisa_a\[6\] VGND sg13g2_inv_1
XFILLER_118_558 VPWR VGND sg13g2_fill_1
XFILLER_66_0 VPWR VGND sg13g2_decap_8
XFILLER_118_569 VPWR VGND sg13g2_decap_8
XFILLER_106_709 VPWR VGND sg13g2_fill_2
XFILLER_105_208 VPWR VGND sg13g2_fill_1
XFILLER_114_797 VPWR VGND sg13g2_decap_8
Xfanout105 net106 net105 VPWR VGND sg13g2_buf_2
XFILLER_113_274 VPWR VGND sg13g2_fill_2
XFILLER_102_937 VPWR VGND sg13g2_decap_8
XFILLER_99_497 VPWR VGND sg13g2_fill_2
Xfanout138 net139 net138 VPWR VGND sg13g2_buf_2
Xfanout116 net119 net116 VPWR VGND sg13g2_buf_2
Xfanout127 net128 net127 VPWR VGND sg13g2_buf_2
XFILLER_59_328 VPWR VGND sg13g2_fill_2
XFILLER_101_447 VPWR VGND sg13g2_decap_8
XFILLER_87_659 VPWR VGND sg13g2_decap_8
X_07984_ _02255_ fp16_sum_pipe.exp_mant_logic0.a\[10\] _02250_ fp16_sum_pipe.seg_reg0.q\[25\]
+ net1775 VPWR VGND sg13g2_a22oi_1
X_09723_ _03839_ _03828_ acc_sum.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_103_13 VPWR VGND sg13g2_fill_1
X_09654_ _03771_ _03728_ _03726_ VPWR VGND sg13g2_nand2_1
XFILLER_95_692 VPWR VGND sg13g2_fill_2
XFILLER_83_832 VPWR VGND sg13g2_fill_1
XFILLER_28_726 VPWR VGND sg13g2_decap_4
XFILLER_103_57 VPWR VGND sg13g2_fill_2
XFILLER_103_46 VPWR VGND sg13g2_decap_8
XFILLER_94_191 VPWR VGND sg13g2_decap_8
X_08605_ _02827_ VPWR _02828_ VGND _02774_ _02826_ sg13g2_o21ai_1
XFILLER_83_876 VPWR VGND sg13g2_fill_1
XFILLER_82_353 VPWR VGND sg13g2_decap_8
XFILLER_43_718 VPWR VGND sg13g2_decap_8
XFILLER_103_79 VPWR VGND sg13g2_fill_2
X_09585_ _03702_ _02806_ _03673_ VPWR VGND sg13g2_nand2_1
XFILLER_27_269 VPWR VGND sg13g2_decap_8
X_08536_ _02760_ acc_sum.op_sign_logic0.mantisa_a\[1\] VPWR VGND acc_sum.op_sign_logic0.mantisa_b\[1\]
+ sg13g2_nand2b_2
XFILLER_36_792 VPWR VGND sg13g2_fill_2
XFILLER_24_932 VPWR VGND sg13g2_decap_8
X_08467_ _02699_ net1647 _02698_ VPWR VGND sg13g2_nand2_1
XFILLER_51_784 VPWR VGND sg13g2_decap_8
XFILLER_23_464 VPWR VGND sg13g2_fill_1
X_07418_ _01754_ net1890 acc\[0\] VPWR VGND sg13g2_nand2_1
X_08398_ VGND VPWR _02592_ _02629_ _02635_ _02634_ sg13g2_a21oi_1
X_07349_ _01708_ VPWR _01476_ VGND acc_sub.reg2en.q\[0\] _01707_ sg13g2_o21ai_1
XFILLER_7_619 VPWR VGND sg13g2_decap_8
XFILLER_12_21 VPWR VGND sg13g2_decap_8
X_10360_ _04403_ _04409_ _04410_ VPWR VGND sg13g2_nor2_1
X_09019_ VGND VPWR _03202_ _03173_ _03205_ _03204_ sg13g2_a21oi_1
XFILLER_105_720 VPWR VGND sg13g2_decap_8
XFILLER_88_36 VPWR VGND sg13g2_decap_8
XFILLER_88_25 VPWR VGND sg13g2_fill_2
XFILLER_3_847 VPWR VGND sg13g2_decap_8
XFILLER_2_302 VPWR VGND sg13g2_fill_2
X_10291_ _01192_ _04358_ _04359_ VPWR VGND sg13g2_nand2_1
XFILLER_12_98 VPWR VGND sg13g2_decap_8
XFILLER_105_742 VPWR VGND sg13g2_fill_2
XFILLER_105_731 VPWR VGND sg13g2_decap_8
X_12030_ VPWR _05877_ fpmul.seg_reg0.q\[16\] VGND sg13g2_inv_1
XFILLER_2_346 VPWR VGND sg13g2_decap_8
XFILLER_104_263 VPWR VGND sg13g2_decap_8
XFILLER_104_241 VPWR VGND sg13g2_decap_8
XFILLER_78_659 VPWR VGND sg13g2_decap_4
XFILLER_77_114 VPWR VGND sg13g2_fill_2
XFILLER_120_778 VPWR VGND sg13g2_decap_8
XFILLER_77_169 VPWR VGND sg13g2_decap_8
XFILLER_59_884 VPWR VGND sg13g2_decap_8
XFILLER_59_851 VPWR VGND sg13g2_fill_2
X_13981_ VPWR _00532_ net12 VGND sg13g2_inv_1
XFILLER_100_480 VPWR VGND sg13g2_decap_8
XFILLER_92_128 VPWR VGND sg13g2_fill_2
X_12932_ VGND VPWR net1936 add_result\[3\] _06705_ net1950 sg13g2_a21oi_1
XFILLER_18_214 VPWR VGND sg13g2_fill_1
XFILLER_100_491 VPWR VGND sg13g2_fill_1
XFILLER_85_191 VPWR VGND sg13g2_decap_8
XFILLER_73_342 VPWR VGND sg13g2_fill_2
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_74_898 VPWR VGND sg13g2_fill_1
XFILLER_74_887 VPWR VGND sg13g2_decap_8
X_12863_ _06642_ _06641_ VPWR VGND _06640_ sg13g2_nand2b_2
X_14602_ _00403_ VGND VPWR _01134_ fp16_res_pipe.y\[13\] clknet_leaf_129_clk sg13g2_dfrbpq_2
XFILLER_15_910 VPWR VGND sg13g2_decap_8
X_11814_ net1837 _05714_ _05709_ _05715_ VPWR VGND sg13g2_nand3_1
XFILLER_14_420 VPWR VGND sg13g2_decap_8
XFILLER_18_1004 VPWR VGND sg13g2_decap_8
X_14533_ _00334_ VGND VPWR _01069_ fpdiv.div_out\[8\] clknet_leaf_76_clk sg13g2_dfrbpq_2
X_11745_ _05647_ _05648_ _05646_ _05649_ VPWR VGND sg13g2_nand3_1
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_30_913 VPWR VGND sg13g2_decap_8
XFILLER_105_1007 VPWR VGND sg13g2_decap_8
X_14464_ _00265_ VGND VPWR _01003_ fpmul.seg_reg0.q\[49\] clknet_leaf_93_clk sg13g2_dfrbpq_1
X_13415_ _07086_ VPWR _00796_ VGND _07040_ net1722 sg13g2_o21ai_1
X_11676_ _05580_ _05579_ fp16_sum_pipe.add_renorm0.exp\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_127_322 VPWR VGND sg13g2_decap_8
X_14395_ _00196_ VGND VPWR _00934_ div_result\[8\] clknet_leaf_87_clk sg13g2_dfrbpq_1
X_10627_ VGND VPWR _03565_ _03572_ _04640_ _04633_ sg13g2_a21oi_1
Xplace1808 acc_sum.exp_mant_logic0.a\[6\] net1808 VPWR VGND sg13g2_buf_2
X_13346_ _07047_ _07027_ fp16_res_pipe.x2\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_5_140 VPWR VGND sg13g2_decap_8
X_10558_ _04590_ VPWR _01156_ VGND net1845 _04589_ sg13g2_o21ai_1
XFILLER_127_399 VPWR VGND sg13g2_decap_8
X_13277_ _06993_ _06994_ _06992_ _06995_ VPWR VGND sg13g2_nand3_1
Xplace1819 acc_sum.reg2en.q\[0\] net1819 VPWR VGND sg13g2_buf_1
XFILLER_6_696 VPWR VGND sg13g2_decap_4
X_12228_ _06074_ _05967_ _06073_ VPWR VGND sg13g2_xnor2_1
X_10489_ net1847 fp16_sum_pipe.add_renorm0.mantisa\[8\] _04535_ VPWR VGND sg13g2_nor2_1
XFILLER_111_701 VPWR VGND sg13g2_decap_8
XFILLER_97_935 VPWR VGND sg13g2_decap_8
XFILLER_96_412 VPWR VGND sg13g2_decap_8
XFILLER_69_615 VPWR VGND sg13g2_fill_1
X_12159_ _06003_ _06004_ _05986_ _06005_ VPWR VGND sg13g2_nand3_1
XFILLER_2_891 VPWR VGND sg13g2_decap_8
XFILLER_25_1008 VPWR VGND sg13g2_decap_4
XFILLER_111_789 VPWR VGND sg13g2_decap_8
XFILLER_68_147 VPWR VGND sg13g2_decap_8
XFILLER_110_288 VPWR VGND sg13g2_decap_8
XFILLER_83_117 VPWR VGND sg13g2_decap_8
XFILLER_65_843 VPWR VGND sg13g2_decap_4
XFILLER_65_810 VPWR VGND sg13g2_decap_4
X_09370_ _03519_ VPWR _03520_ VGND _03500_ _03515_ sg13g2_o21ai_1
X_08321_ _02566_ _02565_ VPWR VGND sg13g2_inv_2
XFILLER_60_592 VPWR VGND sg13g2_fill_1
X_08252_ _02501_ _02502_ _02500_ _02503_ VPWR VGND sg13g2_nand3_1
XFILLER_21_924 VPWR VGND sg13g2_decap_8
X_07203_ VPWR _01575_ _01574_ VGND sg13g2_inv_1
XFILLER_119_856 VPWR VGND sg13g2_decap_8
XFILLER_118_300 VPWR VGND sg13g2_decap_4
Xclkbuf_4_12_0_clk clknet_0_clk clknet_4_12_0_clk VPWR VGND sg13g2_buf_8
X_08183_ _02439_ _02440_ _02441_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_489 VPWR VGND sg13g2_fill_1
XFILLER_118_366 VPWR VGND sg13g2_decap_8
X_07134_ acc_sub.op_sign_logic0.mantisa_a\[8\] _01505_ _01506_ VPWR VGND sg13g2_nor2_1
XFILLER_114_572 VPWR VGND sg13g2_decap_8
XFILLER_114_550 VPWR VGND sg13g2_decap_8
XFILLER_0_828 VPWR VGND sg13g2_decap_8
XFILLER_102_756 VPWR VGND sg13g2_decap_8
XFILLER_88_946 VPWR VGND sg13g2_decap_8
XFILLER_87_423 VPWR VGND sg13g2_decap_8
XFILLER_75_618 VPWR VGND sg13g2_decap_4
X_07967_ _02241_ _02234_ _02240_ VPWR VGND sg13g2_nand2_2
XFILLER_114_56 VPWR VGND sg13g2_decap_8
XFILLER_96_990 VPWR VGND sg13g2_decap_8
X_09706_ VGND VPWR _03820_ net1807 _03822_ _03821_ sg13g2_a21oi_1
XFILLER_74_117 VPWR VGND sg13g2_fill_1
XFILLER_68_670 VPWR VGND sg13g2_fill_1
XFILLER_56_821 VPWR VGND sg13g2_decap_4
XFILLER_56_810 VPWR VGND sg13g2_fill_1
X_07898_ _02176_ net1892 acc_sub.x2\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_56_876 VPWR VGND sg13g2_decap_8
XFILLER_55_320 VPWR VGND sg13g2_fill_2
X_09637_ _03754_ _03630_ _03631_ VPWR VGND sg13g2_nand2_1
XFILLER_83_695 VPWR VGND sg13g2_fill_2
XFILLER_55_386 VPWR VGND sg13g2_decap_4
XFILLER_55_364 VPWR VGND sg13g2_fill_2
XFILLER_43_515 VPWR VGND sg13g2_decap_8
XFILLER_15_217 VPWR VGND sg13g2_decap_4
X_09568_ _03685_ _03674_ _03667_ _03684_ _03655_ VPWR VGND sg13g2_a22oi_1
XFILLER_82_183 VPWR VGND sg13g2_decap_4
XFILLER_43_559 VPWR VGND sg13g2_decap_4
X_08519_ _02740_ _02742_ _02743_ VPWR VGND sg13g2_nor2_1
XFILLER_23_250 VPWR VGND sg13g2_fill_1
XFILLER_24_773 VPWR VGND sg13g2_decap_8
X_09499_ _03617_ fp16_res_pipe.exp_mant_logic0.a\[0\] VPWR VGND sg13g2_inv_2
XFILLER_11_401 VPWR VGND sg13g2_fill_2
XFILLER_11_412 VPWR VGND sg13g2_decap_8
XFILLER_12_946 VPWR VGND sg13g2_decap_8
X_11530_ VPWR _05435_ _05434_ VGND sg13g2_inv_1
XFILLER_11_456 VPWR VGND sg13g2_decap_4
XFILLER_23_42 VPWR VGND sg13g2_decap_8
XFILLER_23_294 VPWR VGND sg13g2_decap_8
XFILLER_99_13 VPWR VGND sg13g2_fill_2
X_11461_ VGND VPWR _05382_ net1944 _01046_ _05383_ sg13g2_a21oi_1
X_14180_ VPWR _00731_ net139 VGND sg13g2_inv_1
XFILLER_99_35 VPWR VGND sg13g2_decap_8
X_11392_ _05340_ net1707 fpdiv.div_out\[10\] VPWR VGND sg13g2_nand2_1
X_13200_ _06934_ VPWR _00859_ VGND _06933_ net1713 sg13g2_o21ai_1
XFILLER_20_990 VPWR VGND sg13g2_decap_8
X_10412_ VPWR _04462_ fp16_sum_pipe.reg2en.q\[0\] VGND sg13g2_inv_1
XFILLER_125_837 VPWR VGND sg13g2_decap_8
X_13131_ _06882_ piso.tx_bit_counter\[4\] _00877_ VPWR VGND sg13g2_nor2b_1
X_10343_ VPWR _04393_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[9\] VGND sg13g2_inv_1
XFILLER_124_336 VPWR VGND sg13g2_decap_8
XFILLER_3_622 VPWR VGND sg13g2_fill_1
X_13062_ _05803_ _05805_ _05801_ _06830_ VPWR VGND _05807_ sg13g2_nand4_1
XFILLER_3_688 VPWR VGND sg13g2_decap_4
XFILLER_2_154 VPWR VGND sg13g2_decap_8
X_10274_ _04343_ VPWR _04344_ VGND _04322_ _04124_ sg13g2_o21ai_1
XFILLER_78_423 VPWR VGND sg13g2_decap_8
X_12013_ net1878 _05852_ _05865_ VPWR VGND _05864_ sg13g2_nand3b_1
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_19_556 VPWR VGND sg13g2_decap_8
X_13964_ VPWR _00515_ net18 VGND sg13g2_inv_1
X_12915_ _06689_ VPWR _06690_ VGND net1962 _06687_ sg13g2_o21ai_1
XFILLER_62_802 VPWR VGND sg13g2_decap_4
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_19_589 VPWR VGND sg13g2_decap_8
X_13895_ VPWR _00446_ net11 VGND sg13g2_inv_1
X_12846_ _00016_ net1730 net1701 _06626_ VPWR VGND sg13g2_nand3_1
XFILLER_61_334 VPWR VGND sg13g2_decap_8
XFILLER_34_537 VPWR VGND sg13g2_fill_2
XFILLER_15_773 VPWR VGND sg13g2_decap_8
X_14516_ _00317_ VGND VPWR _01052_ fpdiv.reg_a_out\[7\] clknet_leaf_56_clk sg13g2_dfrbpq_2
X_12777_ VGND VPWR net1958 fpmul.reg_p_out\[15\] _06562_ _06561_ sg13g2_a21oi_1
XFILLER_42_592 VPWR VGND sg13g2_decap_8
XFILLER_14_250 VPWR VGND sg13g2_fill_1
XFILLER_14_283 VPWR VGND sg13g2_decap_8
XFILLER_9_77 VPWR VGND sg13g2_decap_8
X_11728_ _05483_ _05486_ _05632_ VPWR VGND sg13g2_nor2_1
XFILLER_119_119 VPWR VGND sg13g2_decap_8
X_14447_ _00248_ VGND VPWR _00986_ fpmul.seg_reg0.q\[32\] clknet_leaf_97_clk sg13g2_dfrbpq_1
X_11659_ _05564_ _05405_ _05417_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_1012 VPWR VGND sg13g2_fill_2
X_14378_ _00179_ VGND VPWR _00919_ fpmul.reg_b_out\[9\] clknet_leaf_125_clk sg13g2_dfrbpq_2
X_13329_ _07035_ VPWR _00831_ VGND _07034_ net1725 sg13g2_o21ai_1
XFILLER_7_972 VPWR VGND sg13g2_decap_8
XFILLER_6_460 VPWR VGND sg13g2_decap_8
XFILLER_127_196 VPWR VGND sg13g2_decap_8
Xplace1649 _01959_ net1649 VPWR VGND sg13g2_buf_2
Xplace1638 _02475_ net1638 VPWR VGND sg13g2_buf_2
XFILLER_115_369 VPWR VGND sg13g2_fill_1
XFILLER_9_1013 VPWR VGND sg13g2_fill_1
X_08870_ acc_sub.add_renorm0.mantisa\[1\] _03029_ _03056_ _03057_ VPWR VGND sg13g2_nor3_1
XFILLER_97_754 VPWR VGND sg13g2_fill_1
XFILLER_97_743 VPWR VGND sg13g2_decap_8
X_07821_ _02116_ _02117_ _02115_ _02118_ VPWR VGND sg13g2_nand3_1
XFILLER_97_765 VPWR VGND sg13g2_decap_8
XFILLER_96_253 VPWR VGND sg13g2_fill_1
XFILLER_96_242 VPWR VGND sg13g2_decap_8
XFILLER_57_607 VPWR VGND sg13g2_decap_8
XFILLER_29_0 VPWR VGND sg13g2_decap_8
XFILLER_84_415 VPWR VGND sg13g2_decap_8
X_07752_ acc_sub.exp_mant_logic0.b\[6\] acc_sub.exp_mant_logic0.b\[5\] acc_sub.exp_mant_logic0.b\[4\]
+ acc_sub.exp_mant_logic0.b\[3\] _02056_ VPWR VGND sg13g2_nor4_1
X_07683_ _01992_ _01987_ _01991_ VPWR VGND sg13g2_nand2_1
XFILLER_93_982 VPWR VGND sg13g2_decap_8
XFILLER_38_876 VPWR VGND sg13g2_decap_8
XFILLER_25_504 VPWR VGND sg13g2_decap_8
XFILLER_80_643 VPWR VGND sg13g2_fill_1
XFILLER_80_621 VPWR VGND sg13g2_decap_4
XFILLER_64_172 VPWR VGND sg13g2_decap_4
XFILLER_52_334 VPWR VGND sg13g2_decap_8
X_09422_ VPWR _03565_ fp16_res_pipe.add_renorm0.mantisa\[1\] VGND sg13g2_inv_1
XFILLER_25_537 VPWR VGND sg13g2_decap_4
XFILLER_80_665 VPWR VGND sg13g2_decap_8
XFILLER_40_507 VPWR VGND sg13g2_decap_8
X_09353_ net1738 _03477_ _03503_ _03504_ VPWR VGND sg13g2_nand3_1
X_08304_ _02551_ net1774 fp16_sum_pipe.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_21_732 VPWR VGND sg13g2_fill_2
X_09284_ _03376_ _03437_ _03438_ VPWR VGND sg13g2_nor2_1
X_08235_ _02486_ _02487_ _02485_ _02488_ VPWR VGND sg13g2_nand3_1
XFILLER_20_253 VPWR VGND sg13g2_decap_8
XFILLER_20_264 VPWR VGND sg13g2_fill_1
XFILLER_119_664 VPWR VGND sg13g2_decap_4
X_08166_ _02425_ fp16_sum_pipe.exp_mant_logic0.a\[6\] _02408_ _02273_ _02332_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_20_297 VPWR VGND sg13g2_decap_8
X_07117_ _01490_ acc_sub.seg_reg1.q\[21\] VPWR VGND sg13g2_inv_2
XFILLER_109_56 VPWR VGND sg13g2_decap_8
XFILLER_107_837 VPWR VGND sg13g2_decap_8
XFILLER_107_826 VPWR VGND sg13g2_fill_2
XFILLER_118_196 VPWR VGND sg13g2_decap_8
XFILLER_106_347 VPWR VGND sg13g2_decap_8
X_08097_ _02362_ fp16_sum_pipe.exp_mant_logic0.a\[5\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[8\]
+ net1776 VPWR VGND sg13g2_a22oi_1
XFILLER_121_306 VPWR VGND sg13g2_fill_1
Xclkload90 clknet_leaf_82_clk clkload90/Y VPWR VGND sg13g2_inv_4
XFILLER_125_77 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_0_669 VPWR VGND sg13g2_fill_2
X_08999_ VPWR _03185_ _03184_ VGND sg13g2_inv_1
XFILLER_102_597 VPWR VGND sg13g2_fill_2
XFILLER_75_415 VPWR VGND sg13g2_decap_8
XFILLER_47_117 VPWR VGND sg13g2_decap_8
XFILLER_18_42 VPWR VGND sg13g2_decap_8
XFILLER_28_320 VPWR VGND sg13g2_decap_8
XFILLER_16_504 VPWR VGND sg13g2_fill_1
X_10961_ _04966_ _04964_ _04965_ _04963_ _04962_ VPWR VGND sg13g2_a22oi_1
X_12700_ _06479_ VPWR _06509_ VGND net1734 _06508_ sg13g2_o21ai_1
XFILLER_70_120 VPWR VGND sg13g2_fill_1
X_13680_ VPWR _00231_ net69 VGND sg13g2_inv_1
XFILLER_43_334 VPWR VGND sg13g2_decap_8
X_12631_ VPWR _06447_ _06446_ VGND sg13g2_inv_1
XFILLER_71_665 VPWR VGND sg13g2_decap_8
XFILLER_44_868 VPWR VGND sg13g2_decap_8
XFILLER_43_367 VPWR VGND sg13g2_decap_8
X_10892_ VPWR _04902_ fp16_res_pipe.y\[12\] VGND sg13g2_inv_1
XFILLER_71_687 VPWR VGND sg13g2_decap_8
XFILLER_70_175 VPWR VGND sg13g2_decap_8
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_12_721 VPWR VGND sg13g2_decap_8
XFILLER_24_581 VPWR VGND sg13g2_fill_1
X_12562_ _05370_ fpdiv.reg_b_out\[7\] _06377_ _06378_ VPWR VGND sg13g2_nor3_1
X_14301_ _00102_ VGND VPWR _00845_ acc\[11\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_12493_ net1871 fpmul.seg_reg0.q\[5\] _06329_ VPWR VGND sg13g2_nor2_1
X_11513_ _05405_ _05417_ _05418_ VPWR VGND sg13g2_nor2_1
X_11444_ VPWR _05372_ fpdiv.divider0.dividend\[10\] VGND sg13g2_inv_1
X_14232_ _00033_ VGND VPWR _00783_ sipo.shift_reg\[13\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_8_769 VPWR VGND sg13g2_fill_1
XFILLER_109_174 VPWR VGND sg13g2_decap_4
XFILLER_50_84 VPWR VGND sg13g2_decap_8
XFILLER_124_133 VPWR VGND sg13g2_decap_8
X_14163_ VPWR _00714_ net101 VGND sg13g2_inv_1
X_11375_ _05326_ _05227_ acc_sum.exp_mant_logic0.b\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_98_507 VPWR VGND sg13g2_decap_8
X_13114_ _06871_ _06787_ _06870_ VPWR VGND sg13g2_xnor2_1
XFILLER_4_986 VPWR VGND sg13g2_decap_8
XFILLER_3_441 VPWR VGND sg13g2_decap_8
X_14094_ VPWR _00645_ net41 VGND sg13g2_inv_1
X_10326_ _04380_ VPWR _01178_ VGND net1921 _04329_ sg13g2_o21ai_1
XFILLER_78_220 VPWR VGND sg13g2_fill_1
X_13045_ VPWR _06813_ _06812_ VGND sg13g2_inv_1
X_10257_ _04328_ _04326_ _04327_ VPWR VGND sg13g2_nand2_1
XFILLER_121_840 VPWR VGND sg13g2_decap_8
XFILLER_22_7 VPWR VGND sg13g2_decap_8
XFILLER_78_275 VPWR VGND sg13g2_fill_1
XFILLER_66_437 VPWR VGND sg13g2_decap_8
X_10188_ fp16_res_pipe.exp_mant_logic0.b\[6\] fp16_res_pipe.exp_mant_logic0.b\[5\]
+ fp16_res_pipe.exp_mant_logic0.b\[4\] fp16_res_pipe.exp_mant_logic0.b\[3\] _04266_
+ VPWR VGND sg13g2_nor4_1
XFILLER_82_919 VPWR VGND sg13g2_decap_8
XFILLER_78_297 VPWR VGND sg13g2_fill_2
XFILLER_19_320 VPWR VGND sg13g2_decap_8
X_13947_ VPWR _00498_ net97 VGND sg13g2_inv_1
XFILLER_74_470 VPWR VGND sg13g2_decap_8
XFILLER_62_632 VPWR VGND sg13g2_decap_8
XFILLER_90_974 VPWR VGND sg13g2_decap_8
XFILLER_62_654 VPWR VGND sg13g2_fill_1
XFILLER_35_879 VPWR VGND sg13g2_fill_2
X_13878_ VPWR _00429_ net53 VGND sg13g2_inv_1
XFILLER_22_507 VPWR VGND sg13g2_decap_8
X_12829_ _06611_ _06610_ net1959 VPWR VGND sg13g2_nand2_1
XFILLER_61_175 VPWR VGND sg13g2_fill_1
XFILLER_34_378 VPWR VGND sg13g2_decap_8
XFILLER_30_562 VPWR VGND sg13g2_fill_1
XFILLER_30_573 VPWR VGND sg13g2_decap_8
X_08020_ VGND VPWR _02285_ _02236_ _02286_ _02200_ sg13g2_a21oi_1
XFILLER_116_612 VPWR VGND sg13g2_fill_2
XFILLER_116_656 VPWR VGND sg13g2_decap_8
XFILLER_115_133 VPWR VGND sg13g2_decap_8
Xfanout7 net15 net7 VPWR VGND sg13g2_buf_2
XFILLER_118_1006 VPWR VGND sg13g2_decap_8
XFILLER_116_667 VPWR VGND sg13g2_fill_1
X_09971_ _04063_ _04056_ fp16_res_pipe.exp_mant_logic0.a\[9\] VPWR VGND sg13g2_nand2_1
X_08922_ _03106_ _03107_ _03105_ _03109_ VPWR VGND _03108_ sg13g2_nand4_1
XFILLER_97_562 VPWR VGND sg13g2_decap_8
X_08853_ _03040_ net1789 acc_sub.add_renorm0.mantisa\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_112_873 VPWR VGND sg13g2_decap_8
X_08784_ _02971_ acc_sub.add_renorm0.mantisa\[6\] _02970_ VPWR VGND sg13g2_xnor2_1
X_07804_ _02102_ _01989_ net1747 VPWR VGND sg13g2_nand2_1
XFILLER_85_779 VPWR VGND sg13g2_decap_8
XFILLER_85_757 VPWR VGND sg13g2_fill_1
XFILLER_84_234 VPWR VGND sg13g2_fill_2
X_07735_ _02041_ net1779 acc_sub.op_sign_logic0.mantisa_a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_53_643 VPWR VGND sg13g2_decap_4
XFILLER_25_323 VPWR VGND sg13g2_decap_8
XFILLER_26_846 VPWR VGND sg13g2_fill_1
XFILLER_111_35 VPWR VGND sg13g2_decap_8
XFILLER_81_985 VPWR VGND sg13g2_decap_8
X_09405_ _03549_ VPWR _03550_ VGND _03404_ _03417_ sg13g2_o21ai_1
XFILLER_25_367 VPWR VGND sg13g2_decap_4
XFILLER_26_879 VPWR VGND sg13g2_fill_1
X_07597_ _01911_ net1686 _01884_ VPWR VGND sg13g2_nand2_1
XFILLER_40_326 VPWR VGND sg13g2_decap_8
X_09336_ VGND VPWR _03449_ _03415_ _03488_ _03487_ sg13g2_a21oi_1
X_09267_ VPWR _03421_ fp16_res_pipe.op_sign_logic0.mantisa_b\[4\] VGND sg13g2_inv_1
XFILLER_21_595 VPWR VGND sg13g2_decap_8
X_08218_ _02473_ VPWR _01372_ VGND fp16_sum_pipe.reg1en.q\[0\] _02457_ sg13g2_o21ai_1
Xclkbuf_leaf_141_clk clknet_5_1__leaf_clk clknet_leaf_141_clk VPWR VGND sg13g2_buf_8
X_09198_ _03355_ acc_sum.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_inv_2
XFILLER_106_100 VPWR VGND sg13g2_decap_8
XFILLER_20_21 VPWR VGND sg13g2_decap_8
XFILLER_122_604 VPWR VGND sg13g2_fill_1
X_11160_ _05024_ _05120_ _05106_ _05129_ VPWR VGND sg13g2_nor3_1
XFILLER_122_648 VPWR VGND sg13g2_fill_2
XFILLER_106_199 VPWR VGND sg13g2_decap_4
X_11091_ _05064_ _05049_ acc_sum.exp_mant_logic0.b\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_0_400 VPWR VGND sg13g2_decap_8
XFILLER_1_934 VPWR VGND sg13g2_decap_8
X_10111_ _01207_ _04193_ _04194_ VPWR VGND sg13g2_nand2_1
XFILLER_121_147 VPWR VGND sg13g2_decap_8
XFILLER_103_862 VPWR VGND sg13g2_decap_8
XFILLER_96_36 VPWR VGND sg13g2_fill_1
XFILLER_88_540 VPWR VGND sg13g2_fill_2
X_10042_ _04130_ _04128_ _04017_ VPWR VGND sg13g2_nand2_1
XFILLER_102_372 VPWR VGND sg13g2_decap_4
XFILLER_49_938 VPWR VGND sg13g2_decap_8
XFILLER_0_477 VPWR VGND sg13g2_decap_8
XFILLER_102_394 VPWR VGND sg13g2_fill_2
XFILLER_102_383 VPWR VGND sg13g2_decap_8
XFILLER_75_245 VPWR VGND sg13g2_decap_8
XFILLER_75_234 VPWR VGND sg13g2_decap_4
XFILLER_48_459 VPWR VGND sg13g2_decap_8
X_14850_ _00651_ VGND VPWR _01374_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[1\] clknet_leaf_114_clk
+ sg13g2_dfrbpq_2
XFILLER_29_63 VPWR VGND sg13g2_decap_8
X_14781_ _00582_ VGND VPWR _01305_ acc_sub.y\[10\] clknet_5_21__leaf_clk sg13g2_dfrbpq_1
XFILLER_91_716 VPWR VGND sg13g2_fill_2
XFILLER_91_705 VPWR VGND sg13g2_decap_8
X_13801_ VPWR _00352_ net73 VGND sg13g2_inv_1
XFILLER_17_802 VPWR VGND sg13g2_fill_1
X_11993_ _05834_ _05833_ _05846_ _05847_ VPWR VGND sg13g2_a21o_1
X_13732_ VPWR _00283_ net63 VGND sg13g2_inv_1
XFILLER_17_824 VPWR VGND sg13g2_decap_8
XFILLER_72_963 VPWR VGND sg13g2_fill_1
X_10944_ _04950_ VPWR _01130_ VGND fp16_res_pipe.reg3en.q\[0\] _04940_ sg13g2_o21ai_1
XFILLER_16_345 VPWR VGND sg13g2_decap_8
XFILLER_71_462 VPWR VGND sg13g2_decap_8
X_13663_ VPWR _00214_ net36 VGND sg13g2_inv_1
XFILLER_45_84 VPWR VGND sg13g2_decap_8
X_10875_ VGND VPWR _04885_ _04819_ _04886_ _04774_ sg13g2_a21oi_1
X_12614_ VGND VPWR _06421_ fpdiv.div_out\[0\] _06430_ fpdiv.div_out\[1\] sg13g2_a21oi_1
X_13594_ VPWR _00145_ net110 VGND sg13g2_inv_1
XFILLER_31_348 VPWR VGND sg13g2_fill_1
XFILLER_31_359 VPWR VGND sg13g2_decap_8
X_12545_ fpdiv.divider0.divisor\[10\] fpdiv.divider0.divisor\[9\] fpdiv.divider0.divisor\[8\]
+ fpdiv.divider0.divisor\[7\] _06362_ VPWR VGND sg13g2_nor4_1
XFILLER_84_9 VPWR VGND sg13g2_fill_1
XFILLER_8_511 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_132_clk clknet_5_2__leaf_clk clknet_leaf_132_clk VPWR VGND sg13g2_buf_8
X_12476_ VGND VPWR _06250_ _06151_ _06316_ _06135_ sg13g2_a21oi_1
XFILLER_8_566 VPWR VGND sg13g2_decap_8
XFILLER_126_932 VPWR VGND sg13g2_decap_8
XFILLER_125_431 VPWR VGND sg13g2_fill_1
X_14215_ VPWR _00766_ net133 VGND sg13g2_inv_1
X_11427_ VPWR _05361_ fpdiv.reg_a_out\[12\] VGND sg13g2_inv_1
XFILLER_6_56 VPWR VGND sg13g2_decap_8
XFILLER_125_453 VPWR VGND sg13g2_decap_4
X_14146_ VPWR _00697_ net130 VGND sg13g2_inv_1
X_11358_ _05309_ VPWR _05310_ VGND _03357_ _05222_ sg13g2_o21ai_1
XFILLER_4_761 VPWR VGND sg13g2_decap_4
X_10309_ _04372_ net1914 fp16_res_pipe.x2\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_4_783 VPWR VGND sg13g2_decap_8
XFILLER_3_271 VPWR VGND sg13g2_decap_4
XFILLER_113_659 VPWR VGND sg13g2_fill_1
XFILLER_98_359 VPWR VGND sg13g2_decap_8
X_14077_ VPWR _00628_ net137 VGND sg13g2_inv_1
X_11289_ _03339_ _03341_ _03337_ _05249_ VPWR VGND _03343_ sg13g2_nand4_1
XFILLER_112_169 VPWR VGND sg13g2_decap_8
X_13028_ VPWR _06796_ _06795_ VGND sg13g2_inv_1
XFILLER_67_768 VPWR VGND sg13g2_decap_4
XFILLER_81_226 VPWR VGND sg13g2_fill_2
XFILLER_81_215 VPWR VGND sg13g2_decap_8
XFILLER_75_790 VPWR VGND sg13g2_decap_8
XFILLER_63_941 VPWR VGND sg13g2_decap_8
XFILLER_35_632 VPWR VGND sg13g2_decap_8
XFILLER_19_161 VPWR VGND sg13g2_fill_2
XFILLER_81_259 VPWR VGND sg13g2_fill_1
XFILLER_63_974 VPWR VGND sg13g2_decap_8
X_07451_ _01776_ acc_sub.exp_mant_logic0.b\[15\] VPWR VGND sg13g2_inv_2
XFILLER_50_624 VPWR VGND sg13g2_decap_4
XFILLER_22_304 VPWR VGND sg13g2_fill_1
XFILLER_96_0 VPWR VGND sg13g2_fill_2
X_07382_ _01730_ net1886 acc\[12\] VPWR VGND sg13g2_nand2_1
X_09121_ VGND VPWR _03227_ acc_sub.add_renorm0.exp\[1\] _03302_ _03222_ sg13g2_a21oi_1
XFILLER_50_679 VPWR VGND sg13g2_fill_2
XFILLER_31_882 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_123_clk clknet_5_3__leaf_clk clknet_leaf_123_clk VPWR VGND sg13g2_buf_8
XFILLER_31_893 VPWR VGND sg13g2_decap_8
XFILLER_117_921 VPWR VGND sg13g2_decap_8
X_09052_ net1791 acc_sub.add_renorm0.exp\[6\] _03238_ VPWR VGND sg13g2_nor2_1
X_08003_ _02270_ fp16_sum_pipe.exp_mant_logic0.a\[0\] VPWR VGND sg13g2_inv_2
XFILLER_117_998 VPWR VGND sg13g2_decap_8
XFILLER_104_626 VPWR VGND sg13g2_fill_2
XFILLER_104_615 VPWR VGND sg13g2_decap_8
XFILLER_104_659 VPWR VGND sg13g2_decap_8
XFILLER_103_136 VPWR VGND sg13g2_decap_4
X_09954_ _04049_ VPWR _01219_ VGND _04032_ net1831 sg13g2_o21ai_1
X_08905_ VPWR _03092_ _02967_ VGND sg13g2_inv_1
X_09885_ fp16_res_pipe.op_sign_logic0.s_a fp16_res_pipe.exp_mant_logic0.a\[15\] net1831
+ _01223_ VPWR VGND sg13g2_mux2_1
X_08836_ _03022_ VPWR _03023_ VGND net1789 acc_sub.add_renorm0.mantisa\[4\] sg13g2_o21ai_1
XFILLER_66_28 VPWR VGND sg13g2_decap_8
XFILLER_100_887 VPWR VGND sg13g2_decap_4
XFILLER_122_56 VPWR VGND sg13g2_decap_8
X_08767_ _02958_ acc\[3\] net1897 VPWR VGND sg13g2_nand2_1
XFILLER_54_941 VPWR VGND sg13g2_decap_8
XFILLER_38_492 VPWR VGND sg13g2_fill_2
XFILLER_38_481 VPWR VGND sg13g2_decap_8
X_08698_ net1817 acc_sum.add_renorm0.mantisa\[2\] _02912_ VPWR VGND sg13g2_nor2_1
X_07718_ _02025_ _01959_ acc_sub.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_14_805 VPWR VGND sg13g2_decap_8
XFILLER_82_49 VPWR VGND sg13g2_decap_4
XFILLER_81_793 VPWR VGND sg13g2_decap_8
XFILLER_15_21 VPWR VGND sg13g2_decap_8
XFILLER_25_175 VPWR VGND sg13g2_decap_8
XFILLER_26_676 VPWR VGND sg13g2_decap_8
XFILLER_41_646 VPWR VGND sg13g2_decap_8
XFILLER_40_112 VPWR VGND sg13g2_decap_8
XFILLER_51_1004 VPWR VGND sg13g2_decap_8
X_09319_ _03471_ VPWR _03472_ VGND _03384_ _03386_ sg13g2_o21ai_1
XFILLER_40_189 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_114_clk clknet_5_8__leaf_clk clknet_leaf_114_clk VPWR VGND sg13g2_buf_8
X_10591_ _04608_ VPWR _01141_ VGND net1927 _02261_ sg13g2_o21ai_1
XFILLER_127_729 VPWR VGND sg13g2_decap_8
XFILLER_126_217 VPWR VGND sg13g2_decap_8
X_12330_ _06175_ _06169_ _06176_ VPWR VGND sg13g2_nor2b_1
XFILLER_31_42 VPWR VGND sg13g2_decap_8
X_12261_ _06107_ _06106_ _06088_ VPWR VGND sg13g2_nand2b_1
XFILLER_108_965 VPWR VGND sg13g2_decap_8
X_11212_ _05174_ _05175_ _05177_ _05178_ VPWR VGND sg13g2_nor3_1
X_14000_ VPWR _00551_ net13 VGND sg13g2_inv_1
XFILLER_123_946 VPWR VGND sg13g2_decap_8
XFILLER_122_423 VPWR VGND sg13g2_decap_8
XFILLER_107_486 VPWR VGND sg13g2_decap_8
X_12192_ _06038_ _06029_ _06035_ VPWR VGND sg13g2_xnor2_1
XFILLER_122_456 VPWR VGND sg13g2_decap_8
X_11143_ VGND VPWR _05079_ _05031_ _05113_ _05015_ sg13g2_a21oi_1
XFILLER_1_731 VPWR VGND sg13g2_fill_1
X_14902_ _00703_ VGND VPWR _01422_ acc_sub.op_sign_logic0.mantisa_a\[1\] clknet_leaf_61_clk
+ sg13g2_dfrbpq_2
XFILLER_0_285 VPWR VGND sg13g2_decap_8
X_10025_ _04112_ VPWR _04113_ VGND _04036_ net1689 sg13g2_o21ai_1
XFILLER_64_727 VPWR VGND sg13g2_fill_2
XFILLER_48_267 VPWR VGND sg13g2_fill_1
X_14833_ _00634_ VGND VPWR _01357_ fpdiv.divider0.remainder_reg\[12\] clknet_leaf_71_clk
+ sg13g2_dfrbpq_1
XFILLER_63_237 VPWR VGND sg13g2_decap_4
XFILLER_36_429 VPWR VGND sg13g2_decap_8
XFILLER_29_481 VPWR VGND sg13g2_decap_8
XFILLER_91_579 VPWR VGND sg13g2_decap_8
X_14764_ _00565_ VGND VPWR _01288_ acc_sum.exp_mant_logic0.b\[9\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_11976_ VPWR _05830_ _05829_ VGND sg13g2_inv_1
XFILLER_45_974 VPWR VGND sg13g2_decap_8
XFILLER_16_131 VPWR VGND sg13g2_decap_8
X_13715_ VPWR _00266_ net54 VGND sg13g2_inv_1
XFILLER_44_473 VPWR VGND sg13g2_decap_8
X_14695_ _00496_ VGND VPWR _01223_ fp16_res_pipe.op_sign_logic0.s_a clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_10927_ _04743_ VPWR _04935_ VGND _04934_ _04888_ sg13g2_o21ai_1
XFILLER_32_624 VPWR VGND sg13g2_decap_8
X_13646_ VPWR _00197_ net110 VGND sg13g2_inv_1
XFILLER_16_197 VPWR VGND sg13g2_decap_4
XFILLER_60_988 VPWR VGND sg13g2_decap_8
X_10858_ _04870_ _04867_ _04869_ VPWR VGND sg13g2_nand2_1
XFILLER_31_156 VPWR VGND sg13g2_decap_4
XFILLER_32_679 VPWR VGND sg13g2_decap_8
X_13577_ VPWR _00128_ net22 VGND sg13g2_inv_1
Xclkbuf_leaf_105_clk clknet_5_14__leaf_clk clknet_leaf_105_clk VPWR VGND sg13g2_buf_8
X_10789_ fp16_res_pipe.add_renorm0.exp\[3\] net1709 _04801_ VPWR VGND sg13g2_nor2_1
XFILLER_117_217 VPWR VGND sg13g2_decap_8
Xclkbuf_5_17__f_clk clknet_4_8_0_clk clknet_5_17__leaf_clk VPWR VGND sg13g2_buf_8
X_12528_ _06350_ acc_sub.x2\[3\] net1956 VPWR VGND sg13g2_nand2_1
XFILLER_8_341 VPWR VGND sg13g2_decap_8
XFILLER_9_864 VPWR VGND sg13g2_decap_8
X_12459_ _06251_ _06265_ _06148_ _06302_ VPWR VGND sg13g2_nand3_1
XFILLER_114_902 VPWR VGND sg13g2_decap_8
XFILLER_113_401 VPWR VGND sg13g2_decap_8
XFILLER_125_294 VPWR VGND sg13g2_decap_8
XFILLER_114_979 VPWR VGND sg13g2_decap_8
XFILLER_98_123 VPWR VGND sg13g2_fill_1
X_14129_ VPWR _00680_ net117 VGND sg13g2_inv_1
XFILLER_86_318 VPWR VGND sg13g2_decap_8
X_09670_ _03787_ _03782_ acc_sum.y\[15\] VPWR VGND sg13g2_nand2_1
X_08621_ _02841_ _02842_ _02816_ _02840_ _02843_ VPWR VGND sg13g2_nor4_1
XFILLER_39_245 VPWR VGND sg13g2_decap_4
XFILLER_11_0 VPWR VGND sg13g2_decap_8
XFILLER_27_407 VPWR VGND sg13g2_fill_1
XFILLER_82_535 VPWR VGND sg13g2_decap_8
XFILLER_55_749 VPWR VGND sg13g2_decap_8
XFILLER_27_429 VPWR VGND sg13g2_decap_8
X_08552_ VPWR _02776_ acc_sum.op_sign_logic0.mantisa_a\[5\] VGND sg13g2_inv_1
XFILLER_36_941 VPWR VGND sg13g2_decap_8
X_07503_ VPWR _01825_ acc_sub.exp_mant_logic0.b\[8\] VGND sg13g2_inv_1
X_08483_ _02692_ VPWR _02712_ VGND _02667_ _02711_ sg13g2_o21ai_1
XFILLER_51_900 VPWR VGND sg13g2_decap_8
X_07434_ VPWR _01766_ fpdiv.divider0.divisor\[8\] VGND sg13g2_inv_1
XFILLER_62_270 VPWR VGND sg13g2_fill_1
XFILLER_22_101 VPWR VGND sg13g2_decap_8
XFILLER_11_819 VPWR VGND sg13g2_fill_1
XFILLER_22_167 VPWR VGND sg13g2_fill_1
X_07365_ VPWR _01719_ acc_sub.add_renorm0.exp\[2\] VGND sg13g2_inv_1
X_09104_ VGND VPWR _03175_ net1704 _03286_ _03206_ sg13g2_a21oi_1
X_07296_ _01663_ net1744 _01662_ acc_sub.add_renorm0.mantisa\[7\] net1784 VPWR VGND
+ sg13g2_a22oi_1
X_09035_ net1790 _01719_ _03221_ VPWR VGND sg13g2_nor2_1
XFILLER_105_902 VPWR VGND sg13g2_decap_8
XFILLER_117_795 VPWR VGND sg13g2_decap_8
XFILLER_116_250 VPWR VGND sg13g2_decap_8
XFILLER_89_112 VPWR VGND sg13g2_fill_2
XFILLER_2_528 VPWR VGND sg13g2_decap_8
XFILLER_117_56 VPWR VGND sg13g2_decap_8
XFILLER_105_979 VPWR VGND sg13g2_decap_8
X_09937_ VPWR _04033_ _04020_ VGND sg13g2_inv_1
XFILLER_86_841 VPWR VGND sg13g2_decap_8
X_09868_ _03974_ _03684_ _03674_ VPWR VGND sg13g2_nand2_1
XFILLER_19_908 VPWR VGND sg13g2_decap_8
X_08819_ VPWR _03006_ _03004_ VGND sg13g2_inv_1
X_09799_ VGND VPWR _03871_ _03908_ _03913_ _03906_ sg13g2_a21oi_1
XFILLER_100_684 VPWR VGND sg13g2_decap_8
XFILLER_86_896 VPWR VGND sg13g2_fill_1
XFILLER_45_204 VPWR VGND sg13g2_decap_8
X_11830_ _05730_ net1756 add_result\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_26_42 VPWR VGND sg13g2_decap_8
X_11761_ _05663_ _05664_ _05665_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_974 VPWR VGND sg13g2_decap_8
X_13500_ VPWR _00051_ net34 VGND sg13g2_inv_1
XFILLER_41_421 VPWR VGND sg13g2_fill_1
XFILLER_14_646 VPWR VGND sg13g2_decap_4
X_14480_ _00281_ VGND VPWR _01018_ add_result\[5\] clknet_leaf_107_clk sg13g2_dfrbpq_1
XFILLER_41_465 VPWR VGND sg13g2_decap_8
XFILLER_9_105 VPWR VGND sg13g2_decap_8
X_11692_ _05595_ VPWR _05596_ VGND _04591_ _05583_ sg13g2_o21ai_1
X_13431_ _07094_ VPWR _00788_ VGND _07014_ net1719 sg13g2_o21ai_1
X_10643_ VPWR _04656_ fp16_res_pipe.add_renorm0.mantisa\[9\] VGND sg13g2_inv_1
X_13362_ _07055_ _02588_ _06960_ VPWR VGND sg13g2_nand2_2
X_10574_ _04600_ acc_sub.x2\[12\] net1924 VPWR VGND sg13g2_nand2_1
XFILLER_42_63 VPWR VGND sg13g2_decap_8
XFILLER_10_863 VPWR VGND sg13g2_decap_8
XFILLER_127_548 VPWR VGND sg13g2_decap_8
X_12313_ _06159_ net1855 net1869 VPWR VGND sg13g2_nand2_1
XFILLER_5_322 VPWR VGND sg13g2_decap_8
X_13293_ _07006_ _06952_ _07007_ VPWR VGND sg13g2_nor2_1
XFILLER_6_878 VPWR VGND sg13g2_decap_8
XFILLER_123_710 VPWR VGND sg13g2_fill_2
XFILLER_108_784 VPWR VGND sg13g2_fill_1
XFILLER_107_272 VPWR VGND sg13g2_decap_8
X_12244_ _05959_ _06064_ _06090_ VPWR VGND sg13g2_nor2_1
XFILLER_123_743 VPWR VGND sg13g2_decap_8
XFILLER_122_231 VPWR VGND sg13g2_decap_8
XFILLER_107_294 VPWR VGND sg13g2_decap_8
XFILLER_96_638 VPWR VGND sg13g2_decap_4
XFILLER_95_104 VPWR VGND sg13g2_decap_8
X_11126_ _05034_ net1698 _05096_ VPWR VGND sg13g2_nor2_1
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_110_426 VPWR VGND sg13g2_fill_2
XFILLER_95_126 VPWR VGND sg13g2_decap_8
XFILLER_77_841 VPWR VGND sg13g2_decap_4
XFILLER_110_459 VPWR VGND sg13g2_decap_8
XFILLER_67_93 VPWR VGND sg13g2_fill_2
XFILLER_67_71 VPWR VGND sg13g2_fill_1
X_11057_ _05035_ _05034_ _05011_ VPWR VGND sg13g2_nand2_1
XFILLER_64_502 VPWR VGND sg13g2_decap_4
XFILLER_3_1008 VPWR VGND sg13g2_decap_4
XFILLER_77_896 VPWR VGND sg13g2_fill_1
X_10008_ _04096_ _04093_ _04095_ VPWR VGND sg13g2_nand2_1
X_14816_ _00617_ VGND VPWR _01340_ acc_sum.add_renorm0.mantisa\[5\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_92_866 VPWR VGND sg13g2_decap_8
XFILLER_91_354 VPWR VGND sg13g2_decap_8
XFILLER_18_941 VPWR VGND sg13g2_decap_8
XFILLER_33_911 VPWR VGND sg13g2_decap_8
X_11959_ _05816_ VPWR _00981_ VGND net1884 _05815_ sg13g2_o21ai_1
X_14747_ _00548_ VGND VPWR _01275_ fp16_res_pipe.add_renorm0.mantisa\[10\] clknet_leaf_139_clk
+ sg13g2_dfrbpq_2
XFILLER_32_410 VPWR VGND sg13g2_fill_2
XFILLER_33_988 VPWR VGND sg13g2_decap_8
X_14678_ _00479_ VGND VPWR _01206_ fp16_res_pipe.op_sign_logic0.mantisa_a\[4\] clknet_leaf_143_clk
+ sg13g2_dfrbpq_2
XFILLER_60_796 VPWR VGND sg13g2_decap_8
X_13629_ VPWR _00180_ net50 VGND sg13g2_inv_1
XFILLER_34_1010 VPWR VGND sg13g2_decap_4
XFILLER_32_487 VPWR VGND sg13g2_fill_2
X_07150_ VPWR _01522_ _01521_ VGND sg13g2_inv_1
XFILLER_9_650 VPWR VGND sg13g2_fill_1
XFILLER_9_661 VPWR VGND sg13g2_fill_1
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_8_182 VPWR VGND sg13g2_decap_8
XFILLER_59_0 VPWR VGND sg13g2_decap_8
XFILLER_102_905 VPWR VGND sg13g2_decap_8
XFILLER_114_776 VPWR VGND sg13g2_decap_8
Xfanout106 net107 net106 VPWR VGND sg13g2_buf_2
XFILLER_102_916 VPWR VGND sg13g2_decap_8
XFILLER_101_404 VPWR VGND sg13g2_fill_2
XFILLER_99_476 VPWR VGND sg13g2_decap_8
Xfanout117 net119 net117 VPWR VGND sg13g2_buf_2
Xfanout128 net141 net128 VPWR VGND sg13g2_buf_2
XFILLER_59_307 VPWR VGND sg13g2_decap_8
X_09722_ _03838_ _03837_ VPWR VGND sg13g2_inv_2
Xfanout139 net140 net139 VPWR VGND sg13g2_buf_2
XFILLER_47_19 VPWR VGND sg13g2_decap_8
X_07983_ _02254_ VPWR _01388_ VGND _02194_ _02248_ sg13g2_o21ai_1
XFILLER_86_159 VPWR VGND sg13g2_decap_4
XFILLER_28_705 VPWR VGND sg13g2_decap_8
X_09653_ _03768_ _03769_ _03766_ _03770_ VPWR VGND sg13g2_nand3_1
XFILLER_95_671 VPWR VGND sg13g2_decap_8
XFILLER_82_310 VPWR VGND sg13g2_decap_8
XFILLER_103_25 VPWR VGND sg13g2_decap_8
X_09584_ VPWR _03701_ _03700_ VGND sg13g2_inv_1
XFILLER_94_181 VPWR VGND sg13g2_fill_1
XFILLER_83_866 VPWR VGND sg13g2_fill_2
X_08604_ _02827_ acc_sum.op_sign_logic0.mantisa_a\[4\] acc_sum.op_sign_logic0.mantisa_b\[4\]
+ VPWR VGND sg13g2_nand2_1
X_08535_ _02757_ _02758_ _02759_ VPWR VGND sg13g2_nor2_1
XFILLER_42_207 VPWR VGND sg13g2_fill_2
XFILLER_24_911 VPWR VGND sg13g2_decap_8
XFILLER_35_281 VPWR VGND sg13g2_fill_1
XFILLER_23_421 VPWR VGND sg13g2_fill_2
X_08466_ _02698_ _02675_ _02674_ VPWR VGND sg13g2_xnor2_1
XFILLER_51_763 VPWR VGND sg13g2_decap_8
XFILLER_23_443 VPWR VGND sg13g2_decap_8
XFILLER_24_988 VPWR VGND sg13g2_decap_8
X_07417_ _01753_ acc_sub.exp_mant_logic0.a\[0\] VPWR VGND sg13g2_inv_2
X_08397_ _02633_ _02622_ _02631_ _02634_ VPWR VGND _02624_ sg13g2_nand4_1
XFILLER_11_627 VPWR VGND sg13g2_decap_4
X_07348_ _01708_ _01587_ acc_sub.reg2en.q\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_109_515 VPWR VGND sg13g2_fill_1
XFILLER_10_126 VPWR VGND sg13g2_decap_8
XFILLER_109_548 VPWR VGND sg13g2_fill_1
XFILLER_6_119 VPWR VGND sg13g2_decap_8
X_07279_ _01647_ acc_sub.add_renorm0.mantisa\[8\] VPWR VGND sg13g2_inv_2
XFILLER_109_559 VPWR VGND sg13g2_fill_2
XFILLER_12_77 VPWR VGND sg13g2_decap_8
X_09018_ _03160_ _03203_ _03204_ VPWR VGND sg13g2_nor2_1
XFILLER_3_826 VPWR VGND sg13g2_decap_8
X_10290_ _04359_ net1763 fp16_res_pipe.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_120_757 VPWR VGND sg13g2_decap_8
X_13980_ VPWR _00531_ net13 VGND sg13g2_inv_1
X_12931_ _00009_ net1731 net1702 _06704_ VPWR VGND sg13g2_nand3_1
XFILLER_46_502 VPWR VGND sg13g2_fill_2
XFILLER_73_321 VPWR VGND sg13g2_decap_4
X_12862_ VGND VPWR _04940_ net1910 _06641_ net1923 sg13g2_a21oi_1
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_18_259 VPWR VGND sg13g2_decap_8
XFILLER_46_579 VPWR VGND sg13g2_decap_8
X_11813_ _05714_ _05496_ _05713_ _05710_ _05491_ VPWR VGND sg13g2_a22oi_1
X_14601_ _00402_ VGND VPWR _01133_ fp16_res_pipe.y\[12\] clknet_leaf_129_clk sg13g2_dfrbpq_1
XFILLER_27_771 VPWR VGND sg13g2_fill_2
X_12793_ _06573_ _06577_ _06563_ _00909_ VPWR VGND sg13g2_nand3_1
X_14532_ _00333_ VGND VPWR _01068_ fpdiv.div_out\[7\] clknet_leaf_77_clk sg13g2_dfrbpq_1
XFILLER_41_251 VPWR VGND sg13g2_decap_8
XFILLER_14_465 VPWR VGND sg13g2_fill_2
XFILLER_15_966 VPWR VGND sg13g2_decap_8
X_11744_ _05489_ _05648_ VPWR VGND sg13g2_inv_4
X_14463_ _00264_ VGND VPWR _01002_ fpmul.seg_reg0.q\[48\] clknet_leaf_92_clk sg13g2_dfrbpq_1
XFILLER_42_796 VPWR VGND sg13g2_fill_1
X_11675_ _04585_ _05578_ _05579_ VPWR VGND sg13g2_nor2_1
X_13414_ _07086_ net1722 instr\[10\] VPWR VGND sg13g2_nand2_1
X_10626_ _04639_ _04615_ _04638_ VPWR VGND sg13g2_xnor2_1
XFILLER_30_969 VPWR VGND sg13g2_decap_8
XFILLER_127_301 VPWR VGND sg13g2_decap_8
X_14394_ _00195_ VGND VPWR _00933_ div_result\[7\] clknet_leaf_88_clk sg13g2_dfrbpq_1
XFILLER_115_507 VPWR VGND sg13g2_decap_8
X_13345_ VPWR _07046_ sipo.word\[7\] VGND sg13g2_inv_1
Xplace1809 acc_sum.exp_mant_logic0.a\[5\] net1809 VPWR VGND sg13g2_buf_2
XFILLER_6_642 VPWR VGND sg13g2_decap_4
XFILLER_10_682 VPWR VGND sg13g2_decap_4
X_10557_ _04590_ fp16_sum_pipe.seg_reg0.q\[25\] net1845 VPWR VGND sg13g2_nand2_1
XFILLER_127_378 VPWR VGND sg13g2_decap_8
X_13276_ _06994_ net1743 sipo.word\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_52_7 VPWR VGND sg13g2_decap_8
XFILLER_6_664 VPWR VGND sg13g2_decap_4
X_10488_ _04534_ _04454_ _04533_ VPWR VGND sg13g2_xnor2_1
X_12227_ _06073_ net1858 net1865 VPWR VGND sg13g2_nand2_1
XFILLER_97_914 VPWR VGND sg13g2_decap_8
XFILLER_2_870 VPWR VGND sg13g2_decap_8
XFILLER_123_595 VPWR VGND sg13g2_decap_8
XFILLER_96_446 VPWR VGND sg13g2_decap_8
XFILLER_69_649 VPWR VGND sg13g2_decap_4
X_12158_ _06001_ _05987_ _05999_ _06004_ VPWR VGND sg13g2_nand3_1
XFILLER_1_380 VPWR VGND sg13g2_decap_8
XFILLER_111_768 VPWR VGND sg13g2_decap_8
X_11109_ VPWR _05079_ _05078_ VGND sg13g2_inv_1
X_12089_ VGND VPWR _05903_ net1868 _05935_ _05934_ sg13g2_a21oi_1
XFILLER_110_278 VPWR VGND sg13g2_decap_4
XFILLER_77_682 VPWR VGND sg13g2_fill_1
XFILLER_65_822 VPWR VGND sg13g2_decap_8
XFILLER_37_524 VPWR VGND sg13g2_decap_8
XFILLER_65_866 VPWR VGND sg13g2_fill_2
XFILLER_65_855 VPWR VGND sg13g2_decap_8
XFILLER_94_91 VPWR VGND sg13g2_decap_8
XFILLER_80_836 VPWR VGND sg13g2_decap_8
XFILLER_37_568 VPWR VGND sg13g2_fill_2
XFILLER_18_771 VPWR VGND sg13g2_decap_8
XFILLER_25_719 VPWR VGND sg13g2_decap_8
XFILLER_91_184 VPWR VGND sg13g2_decap_4
X_08320_ _02565_ _02561_ _02564_ VPWR VGND sg13g2_nand2_1
XFILLER_21_903 VPWR VGND sg13g2_decap_8
X_08251_ _02502_ _02343_ net1842 VPWR VGND sg13g2_nand2_1
XFILLER_20_413 VPWR VGND sg13g2_decap_8
X_07202_ _01573_ VPWR _01574_ VGND _01544_ _01571_ sg13g2_o21ai_1
XFILLER_119_835 VPWR VGND sg13g2_decap_8
X_08182_ _02440_ _02378_ fp16_sum_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
X_07133_ VPWR _01505_ acc_sub.op_sign_logic0.mantisa_b\[8\] VGND sg13g2_inv_1
XFILLER_127_890 VPWR VGND sg13g2_decap_8
XFILLER_87_402 VPWR VGND sg13g2_decap_8
XFILLER_0_807 VPWR VGND sg13g2_decap_8
XFILLER_102_735 VPWR VGND sg13g2_decap_8
XFILLER_101_223 VPWR VGND sg13g2_decap_4
XFILLER_101_212 VPWR VGND sg13g2_decap_8
XFILLER_101_234 VPWR VGND sg13g2_fill_2
X_07966_ VPWR VGND _02191_ _02239_ _02237_ _02187_ _02240_ _02184_ sg13g2_a221oi_1
XFILLER_114_35 VPWR VGND sg13g2_decap_8
X_09705_ net1807 acc_sum.add_renorm0.exp\[6\] _03821_ VPWR VGND sg13g2_nor2_1
XFILLER_28_524 VPWR VGND sg13g2_decap_8
X_09636_ _03753_ _03666_ _03652_ VPWR VGND sg13g2_nand2_1
XFILLER_95_490 VPWR VGND sg13g2_fill_2
X_07897_ _02175_ VPWR _01395_ VGND net1891 _02156_ sg13g2_o21ai_1
Xclkbuf_leaf_94_clk clknet_5_13__leaf_clk clknet_leaf_94_clk VPWR VGND sg13g2_buf_8
XFILLER_83_674 VPWR VGND sg13g2_decap_8
XFILLER_83_663 VPWR VGND sg13g2_fill_1
XFILLER_15_207 VPWR VGND sg13g2_fill_1
X_09567_ _03633_ _03660_ _03684_ VPWR VGND sg13g2_nor2_2
XFILLER_24_730 VPWR VGND sg13g2_fill_2
X_08518_ VPWR _02742_ _02741_ VGND sg13g2_inv_1
X_09498_ _03616_ VPWR _01242_ VGND net1916 _03615_ sg13g2_o21ai_1
X_08449_ _02681_ _02682_ _02683_ VPWR VGND sg13g2_nor2_1
XFILLER_12_925 VPWR VGND sg13g2_decap_8
XFILLER_23_21 VPWR VGND sg13g2_decap_8
X_11460_ net1946 fpdiv.divider0.dividend\[5\] _05383_ VPWR VGND sg13g2_nor2_1
X_11391_ _05339_ fpdiv.div_out\[9\] VPWR VGND sg13g2_inv_2
XFILLER_23_98 VPWR VGND sg13g2_fill_1
XFILLER_125_816 VPWR VGND sg13g2_decap_8
XFILLER_124_315 VPWR VGND sg13g2_decap_8
XFILLER_109_378 VPWR VGND sg13g2_fill_1
XFILLER_109_367 VPWR VGND sg13g2_decap_8
XFILLER_3_601 VPWR VGND sg13g2_decap_8
X_10342_ VPWR _04392_ _04391_ VGND sg13g2_inv_1
X_13061_ _05813_ _05819_ _05811_ _06829_ VPWR VGND sg13g2_nand3_1
XFILLER_3_634 VPWR VGND sg13g2_fill_1
X_12012_ _05851_ _05850_ _05864_ VPWR VGND sg13g2_nor2_1
XFILLER_3_667 VPWR VGND sg13g2_decap_8
XFILLER_2_133 VPWR VGND sg13g2_decap_8
X_10273_ _04343_ net1643 fp16_res_pipe.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_120_510 VPWR VGND sg13g2_fill_2
XFILLER_78_413 VPWR VGND sg13g2_fill_1
XFILLER_120_543 VPWR VGND sg13g2_decap_8
XFILLER_78_457 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_19_524 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_85_clk clknet_5_25__leaf_clk clknet_leaf_85_clk VPWR VGND sg13g2_buf_8
XFILLER_58_192 VPWR VGND sg13g2_fill_1
XFILLER_58_181 VPWR VGND sg13g2_decap_8
X_13963_ VPWR _00514_ net18 VGND sg13g2_inv_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_104_90 VPWR VGND sg13g2_fill_1
XFILLER_73_162 VPWR VGND sg13g2_decap_8
X_12914_ _06689_ _06688_ net1961 VPWR VGND sg13g2_nand2_1
X_13894_ VPWR _00445_ net30 VGND sg13g2_inv_1
X_12845_ _06624_ _06625_ _06615_ _00905_ VPWR VGND sg13g2_nand3_1
XFILLER_74_696 VPWR VGND sg13g2_decap_8
XFILLER_73_195 VPWR VGND sg13g2_fill_1
XFILLER_62_858 VPWR VGND sg13g2_decap_8
X_12776_ _06561_ _06559_ VPWR VGND sg13g2_inv_2
XFILLER_62_869 VPWR VGND sg13g2_fill_1
XFILLER_61_357 VPWR VGND sg13g2_fill_1
X_14515_ _00316_ VGND VPWR _01051_ fpdiv.divider0.dividend\[10\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_1
XFILLER_70_891 VPWR VGND sg13g2_fill_2
XFILLER_30_722 VPWR VGND sg13g2_fill_1
X_11727_ VPWR VGND _05496_ net1757 _05630_ _05491_ _05631_ _05614_ sg13g2_a221oi_1
XFILLER_9_56 VPWR VGND sg13g2_decap_8
XFILLER_30_755 VPWR VGND sg13g2_decap_8
XFILLER_80_71 VPWR VGND sg13g2_fill_2
X_14446_ _00247_ VGND VPWR _00985_ fpmul.seg_reg0.q\[31\] clknet_leaf_97_clk sg13g2_dfrbpq_1
X_11658_ VPWR _05563_ _05562_ VGND sg13g2_inv_1
X_14377_ _00178_ VGND VPWR _00918_ fpmul.reg_b_out\[8\] clknet_leaf_125_clk sg13g2_dfrbpq_2
XFILLER_7_951 VPWR VGND sg13g2_decap_8
X_10609_ _04622_ _04621_ net1826 VPWR VGND sg13g2_nand2_1
XFILLER_11_980 VPWR VGND sg13g2_decap_8
X_11589_ VPWR _05494_ _05493_ VGND sg13g2_inv_1
XFILLER_127_175 VPWR VGND sg13g2_decap_8
X_13328_ _07035_ net1725 fp16_res_pipe.x2\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_116_849 VPWR VGND sg13g2_decap_8
Xplace1639 _02352_ net1639 VPWR VGND sg13g2_buf_2
X_13259_ _06981_ acc_sub.y\[12\] net1711 acc_sum.y\[12\] net1728 VPWR VGND sg13g2_a22oi_1
XFILLER_124_893 VPWR VGND sg13g2_decap_8
XFILLER_69_413 VPWR VGND sg13g2_fill_2
X_07820_ _02117_ net1650 acc_sub.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_69_468 VPWR VGND sg13g2_decap_8
XFILLER_69_446 VPWR VGND sg13g2_decap_8
XFILLER_97_788 VPWR VGND sg13g2_decap_8
XFILLER_96_265 VPWR VGND sg13g2_decap_8
X_07751_ acc_sub.exp_mant_logic0.b\[14\] acc_sub.exp_mant_logic0.b\[13\] acc_sub.exp_mant_logic0.b\[12\]
+ acc_sub.exp_mant_logic0.b\[11\] _02055_ VPWR VGND sg13g2_nor4_1
XFILLER_69_479 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_76_clk clknet_5_27__leaf_clk clknet_leaf_76_clk VPWR VGND sg13g2_buf_8
XFILLER_38_855 VPWR VGND sg13g2_fill_2
X_07682_ _01991_ _01989_ _01869_ VPWR VGND sg13g2_nand2_1
XFILLER_93_961 VPWR VGND sg13g2_decap_8
XFILLER_65_652 VPWR VGND sg13g2_decap_8
XFILLER_64_151 VPWR VGND sg13g2_decap_8
XFILLER_52_302 VPWR VGND sg13g2_decap_8
XFILLER_37_387 VPWR VGND sg13g2_decap_8
X_09421_ _03564_ VPWR _01267_ VGND _03560_ _03561_ sg13g2_o21ai_1
X_09352_ _03503_ _03377_ _03476_ VPWR VGND sg13g2_nand2b_1
XFILLER_52_379 VPWR VGND sg13g2_decap_4
X_08303_ _02550_ _02549_ net1638 VPWR VGND sg13g2_nand2_1
XFILLER_21_711 VPWR VGND sg13g2_decap_8
XFILLER_33_571 VPWR VGND sg13g2_fill_2
X_09283_ VPWR _03437_ _03436_ VGND sg13g2_inv_1
XFILLER_21_744 VPWR VGND sg13g2_decap_8
XFILLER_33_593 VPWR VGND sg13g2_decap_8
X_08234_ _02487_ _02343_ _02472_ VPWR VGND sg13g2_nand2_1
XFILLER_21_766 VPWR VGND sg13g2_decap_8
XFILLER_119_643 VPWR VGND sg13g2_decap_8
X_08165_ _02421_ _02423_ _02424_ VPWR VGND sg13g2_nor2_1
XFILLER_118_175 VPWR VGND sg13g2_decap_8
XFILLER_109_35 VPWR VGND sg13g2_decap_8
Xclkload80 clknet_leaf_34_clk clkload80/Y VPWR VGND sg13g2_inv_4
XFILLER_69_39 VPWR VGND sg13g2_decap_8
X_08096_ _02361_ net1639 _02360_ VPWR VGND sg13g2_nand2_1
XFILLER_122_819 VPWR VGND sg13g2_decap_8
Xclkload91 clknet_leaf_88_clk clkload91/Y VPWR VGND sg13g2_inv_4
XFILLER_115_893 VPWR VGND sg13g2_decap_8
XFILLER_114_381 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_125_56 VPWR VGND sg13g2_decap_8
XFILLER_102_543 VPWR VGND sg13g2_fill_2
XFILLER_76_906 VPWR VGND sg13g2_fill_2
X_08998_ _03184_ _01715_ _03140_ VPWR VGND sg13g2_xnor2_1
XFILLER_85_38 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_67_clk clknet_5_31__leaf_clk clknet_leaf_67_clk VPWR VGND sg13g2_buf_8
XFILLER_87_298 VPWR VGND sg13g2_decap_8
XFILLER_75_449 VPWR VGND sg13g2_decap_8
XFILLER_18_21 VPWR VGND sg13g2_decap_8
XFILLER_28_310 VPWR VGND sg13g2_fill_1
X_10960_ VGND VPWR _04744_ _04841_ _04965_ net1771 sg13g2_a21oi_1
XFILLER_29_899 VPWR VGND sg13g2_decap_8
X_09619_ _03736_ _03735_ _03713_ VPWR VGND sg13g2_nand2_1
XFILLER_84_994 VPWR VGND sg13g2_decap_8
XFILLER_83_471 VPWR VGND sg13g2_decap_8
X_10891_ _01134_ _04900_ _04901_ VPWR VGND sg13g2_nand2_1
XFILLER_28_376 VPWR VGND sg13g2_fill_2
X_12630_ VGND VPWR _06421_ fpdiv.div_out\[5\] _06446_ _06445_ sg13g2_a21oi_1
XFILLER_70_187 VPWR VGND sg13g2_decap_8
XFILLER_54_1013 VPWR VGND sg13g2_fill_1
XFILLER_52_891 VPWR VGND sg13g2_decap_8
XFILLER_34_42 VPWR VGND sg13g2_decap_8
XFILLER_24_560 VPWR VGND sg13g2_decap_4
X_12561_ VPWR _06377_ _06376_ VGND sg13g2_inv_1
XFILLER_15_1008 VPWR VGND sg13g2_decap_4
X_14300_ _00101_ VGND VPWR _00844_ acc\[10\] clknet_leaf_48_clk sg13g2_dfrbpq_2
X_12492_ _06328_ _06240_ _06327_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_726 VPWR VGND sg13g2_decap_4
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_12_788 VPWR VGND sg13g2_fill_2
X_11512_ _05417_ _05416_ VPWR VGND _05408_ sg13g2_nand2b_2
XFILLER_126_0 VPWR VGND sg13g2_decap_8
XFILLER_109_120 VPWR VGND sg13g2_decap_4
X_11443_ _05371_ VPWR _01052_ VGND net1944 _05370_ sg13g2_o21ai_1
X_14231_ _00032_ VGND VPWR _00782_ sipo.shift_reg\[12\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_7_247 VPWR VGND sg13g2_decap_8
XFILLER_125_613 VPWR VGND sg13g2_decap_4
XFILLER_109_142 VPWR VGND sg13g2_fill_2
X_14162_ VPWR _00713_ net103 VGND sg13g2_inv_1
XFILLER_50_63 VPWR VGND sg13g2_decap_8
XFILLER_124_112 VPWR VGND sg13g2_decap_8
X_13113_ _06870_ _06869_ _06784_ VPWR VGND sg13g2_nand2_1
X_11374_ _03355_ _05143_ _05325_ VPWR VGND sg13g2_nor2_1
XFILLER_3_420 VPWR VGND sg13g2_decap_8
XFILLER_125_668 VPWR VGND sg13g2_fill_2
XFILLER_106_871 VPWR VGND sg13g2_decap_8
X_14093_ VPWR _00644_ net40 VGND sg13g2_inv_1
XFILLER_4_965 VPWR VGND sg13g2_decap_8
X_10325_ _04380_ net1920 fp16_res_pipe.x2\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_124_189 VPWR VGND sg13g2_decap_8
XFILLER_79_733 VPWR VGND sg13g2_decap_8
X_13044_ _06759_ _06811_ _06812_ VPWR VGND sg13g2_nor2_1
XFILLER_3_497 VPWR VGND sg13g2_decap_8
X_10256_ _04327_ _04190_ net1830 VPWR VGND sg13g2_nand2_1
XFILLER_120_340 VPWR VGND sg13g2_decap_8
XFILLER_78_254 VPWR VGND sg13g2_fill_2
XFILLER_78_243 VPWR VGND sg13g2_decap_8
XFILLER_78_232 VPWR VGND sg13g2_decap_8
XFILLER_59_83 VPWR VGND sg13g2_fill_1
XFILLER_121_896 VPWR VGND sg13g2_decap_8
XFILLER_93_213 VPWR VGND sg13g2_fill_1
XFILLER_66_416 VPWR VGND sg13g2_decap_8
X_10187_ fp16_res_pipe.exp_mant_logic0.b\[14\] fp16_res_pipe.exp_mant_logic0.b\[13\]
+ fp16_res_pipe.exp_mant_logic0.b\[12\] fp16_res_pipe.exp_mant_logic0.b\[11\] _04265_
+ VPWR VGND sg13g2_nor4_1
Xclkbuf_leaf_58_clk clknet_5_30__leaf_clk clknet_leaf_58_clk VPWR VGND sg13g2_buf_8
XFILLER_15_7 VPWR VGND sg13g2_decap_8
Xclkbuf_4_11_0_clk clknet_0_clk clknet_4_11_0_clk VPWR VGND sg13g2_buf_8
XFILLER_75_71 VPWR VGND sg13g2_decap_8
XFILLER_47_663 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
X_13946_ VPWR _00497_ net29 VGND sg13g2_inv_1
XFILLER_19_343 VPWR VGND sg13g2_fill_2
XFILLER_62_611 VPWR VGND sg13g2_decap_8
XFILLER_19_398 VPWR VGND sg13g2_fill_1
XFILLER_90_953 VPWR VGND sg13g2_decap_8
X_13877_ VPWR _00428_ net53 VGND sg13g2_inv_1
XFILLER_34_335 VPWR VGND sg13g2_decap_8
X_12828_ VPWR _06610_ fpmul.reg_p_out\[12\] VGND sg13g2_inv_1
XFILLER_61_154 VPWR VGND sg13g2_decap_8
XFILLER_91_92 VPWR VGND sg13g2_decap_4
XFILLER_91_70 VPWR VGND sg13g2_fill_1
XFILLER_61_198 VPWR VGND sg13g2_decap_8
X_12759_ fpmul.reg_b_out\[1\] fp16_res_pipe.x2\[1\] net1957 _00911_ VPWR VGND sg13g2_mux2_1
XFILLER_15_593 VPWR VGND sg13g2_decap_8
X_14429_ _00230_ VGND VPWR _00968_ fpmul.seg_reg0.q\[14\] clknet_leaf_81_clk sg13g2_dfrbpq_1
XFILLER_115_112 VPWR VGND sg13g2_decap_8
XFILLER_7_781 VPWR VGND sg13g2_decap_4
Xfanout8 net15 net8 VPWR VGND sg13g2_buf_2
XFILLER_116_679 VPWR VGND sg13g2_decap_8
XFILLER_104_819 VPWR VGND sg13g2_decap_8
X_09970_ _04062_ _04052_ fp16_res_pipe.exp_mant_logic0.b\[9\] VPWR VGND sg13g2_nand2_1
X_08921_ _03108_ _03094_ _03001_ VPWR VGND sg13g2_nand2_1
XFILLER_115_189 VPWR VGND sg13g2_decap_8
XFILLER_41_0 VPWR VGND sg13g2_decap_8
XFILLER_112_852 VPWR VGND sg13g2_decap_8
XFILLER_97_541 VPWR VGND sg13g2_decap_8
XFILLER_69_232 VPWR VGND sg13g2_decap_4
X_07803_ _01415_ _02100_ _02101_ VPWR VGND sg13g2_nand2_1
XFILLER_57_416 VPWR VGND sg13g2_fill_2
X_08783_ acc_sub.add_renorm0.mantisa\[5\] acc_sub.add_renorm0.mantisa\[4\] _02969_
+ _02970_ VPWR VGND sg13g2_nand3_1
XFILLER_111_395 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_49_clk clknet_5_22__leaf_clk clknet_leaf_49_clk VPWR VGND sg13g2_buf_8
XFILLER_85_747 VPWR VGND sg13g2_decap_4
X_07734_ _02040_ _02039_ net1641 VPWR VGND sg13g2_nand2_1
XFILLER_66_961 VPWR VGND sg13g2_fill_1
XFILLER_38_652 VPWR VGND sg13g2_decap_4
XFILLER_26_814 VPWR VGND sg13g2_fill_2
X_07665_ net1660 _01974_ _01975_ VPWR VGND sg13g2_nor2b_2
XFILLER_77_1013 VPWR VGND sg13g2_fill_1
XFILLER_38_685 VPWR VGND sg13g2_fill_1
XFILLER_37_184 VPWR VGND sg13g2_fill_2
XFILLER_37_173 VPWR VGND sg13g2_decap_4
XFILLER_111_14 VPWR VGND sg13g2_decap_8
XFILLER_81_964 VPWR VGND sg13g2_decap_8
XFILLER_38_1008 VPWR VGND sg13g2_decap_4
X_09404_ VPWR _03549_ _03406_ VGND sg13g2_inv_1
X_07596_ _01910_ _01909_ _01817_ VPWR VGND sg13g2_nand2_1
XFILLER_80_485 VPWR VGND sg13g2_decap_8
XFILLER_52_198 VPWR VGND sg13g2_fill_1
XFILLER_52_187 VPWR VGND sg13g2_decap_8
XFILLER_34_891 VPWR VGND sg13g2_decap_8
X_09335_ VPWR _03487_ _03413_ VGND sg13g2_inv_1
X_09266_ _03419_ VPWR _03420_ VGND _03408_ _03417_ sg13g2_o21ai_1
X_08217_ net1843 _02472_ _02244_ _02473_ VPWR VGND sg13g2_nand3_1
XFILLER_101_1011 VPWR VGND sg13g2_fill_2
X_09197_ _03354_ VPWR _01281_ VGND net1906 _03353_ sg13g2_o21ai_1
XFILLER_5_707 VPWR VGND sg13g2_decap_8
XFILLER_119_484 VPWR VGND sg13g2_decap_8
XFILLER_4_239 VPWR VGND sg13g2_decap_8
X_08148_ _02305_ _02407_ _02408_ VPWR VGND sg13g2_nor2b_2
XFILLER_107_679 VPWR VGND sg13g2_fill_2
X_08079_ _02345_ _02343_ VPWR VGND sg13g2_inv_2
XFILLER_20_77 VPWR VGND sg13g2_decap_4
XFILLER_122_616 VPWR VGND sg13g2_decap_4
X_11090_ _05063_ VPWR _01097_ VGND _03339_ _05050_ sg13g2_o21ai_1
XFILLER_1_913 VPWR VGND sg13g2_decap_8
XFILLER_20_99 VPWR VGND sg13g2_decap_8
X_10110_ _04194_ fp16_res_pipe.exp_mant_logic0.a\[2\] net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[5\]
+ net1764 VPWR VGND sg13g2_a22oi_1
XFILLER_121_126 VPWR VGND sg13g2_decap_8
XFILLER_103_841 VPWR VGND sg13g2_fill_2
XFILLER_49_917 VPWR VGND sg13g2_decap_8
XFILLER_49_906 VPWR VGND sg13g2_fill_1
XFILLER_102_351 VPWR VGND sg13g2_decap_8
XFILLER_102_340 VPWR VGND sg13g2_decap_4
XFILLER_88_585 VPWR VGND sg13g2_fill_2
XFILLER_0_456 VPWR VGND sg13g2_decap_8
XFILLER_29_42 VPWR VGND sg13g2_decap_8
XFILLER_76_747 VPWR VGND sg13g2_fill_1
XFILLER_75_213 VPWR VGND sg13g2_decap_8
XFILLER_21_1001 VPWR VGND sg13g2_decap_8
X_14780_ _00581_ VGND VPWR _01304_ acc_sub.y\[9\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_13800_ VPWR _00351_ net74 VGND sg13g2_inv_1
X_11992_ _05836_ _05845_ _05846_ VPWR VGND sg13g2_nor2_1
XFILLER_17_814 VPWR VGND sg13g2_fill_1
XFILLER_21_1012 VPWR VGND sg13g2_fill_2
XFILLER_28_140 VPWR VGND sg13g2_decap_8
XFILLER_72_931 VPWR VGND sg13g2_fill_1
XFILLER_72_920 VPWR VGND sg13g2_decap_8
X_13731_ VPWR _00282_ net68 VGND sg13g2_inv_1
XFILLER_16_324 VPWR VGND sg13g2_decap_8
XFILLER_17_847 VPWR VGND sg13g2_fill_2
X_10943_ _04947_ _04949_ _04897_ _04950_ VPWR VGND sg13g2_nand3_1
XFILLER_71_441 VPWR VGND sg13g2_decap_8
XFILLER_45_63 VPWR VGND sg13g2_decap_8
X_13662_ VPWR _00213_ net59 VGND sg13g2_inv_1
XFILLER_44_699 VPWR VGND sg13g2_decap_8
XFILLER_43_176 VPWR VGND sg13g2_decap_8
X_10874_ _04885_ _04884_ _04817_ VPWR VGND sg13g2_nand2_1
X_12613_ _06429_ fpdiv.div_out\[11\] fpdiv.div_out\[2\] VPWR VGND sg13g2_nand2_1
X_13593_ VPWR _00144_ net120 VGND sg13g2_inv_1
XFILLER_43_187 VPWR VGND sg13g2_fill_2
XFILLER_31_327 VPWR VGND sg13g2_decap_8
XFILLER_101_91 VPWR VGND sg13g2_decap_8
X_12544_ fpdiv.divider0.divisor\[6\] fpdiv.divider0.divisor\[5\] fpdiv.divider0.divisor\[4\]
+ fpdiv.reg_b_out\[14\] _06361_ VPWR VGND sg13g2_nor4_1
XFILLER_40_861 VPWR VGND sg13g2_decap_8
XFILLER_61_73 VPWR VGND sg13g2_fill_2
XFILLER_40_894 VPWR VGND sg13g2_decap_8
XFILLER_126_911 VPWR VGND sg13g2_decap_8
X_12475_ _06315_ VPWR _00964_ VGND net1871 _06313_ sg13g2_o21ai_1
X_14214_ VPWR _00765_ net133 VGND sg13g2_inv_1
X_11426_ VGND VPWR _05359_ net1940 _01058_ _05360_ sg13g2_a21oi_1
XFILLER_6_35 VPWR VGND sg13g2_decap_8
XFILLER_126_988 VPWR VGND sg13g2_decap_8
X_14145_ VPWR _00696_ net134 VGND sg13g2_inv_1
X_11357_ _05309_ net1656 acc_sum.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_125_498 VPWR VGND sg13g2_fill_1
XFILLER_113_627 VPWR VGND sg13g2_fill_1
X_14076_ VPWR _00627_ net137 VGND sg13g2_inv_1
X_10308_ _04371_ VPWR _01187_ VGND net1915 _03995_ sg13g2_o21ai_1
XFILLER_98_349 VPWR VGND sg13g2_fill_2
X_13027_ VGND VPWR net1755 fpmul.seg_reg0.q\[6\] _06795_ _06794_ sg13g2_a21oi_1
X_11288_ _03349_ _03355_ _03347_ _05248_ VPWR VGND sg13g2_nand3_1
XFILLER_3_283 VPWR VGND sg13g2_fill_2
XFILLER_94_500 VPWR VGND sg13g2_fill_2
XFILLER_66_202 VPWR VGND sg13g2_fill_2
X_10239_ _04300_ _04140_ _04311_ VPWR VGND sg13g2_nor2_1
XFILLER_121_682 VPWR VGND sg13g2_fill_2
XFILLER_94_544 VPWR VGND sg13g2_fill_1
XFILLER_86_70 VPWR VGND sg13g2_decap_4
XFILLER_67_747 VPWR VGND sg13g2_decap_8
XFILLER_55_909 VPWR VGND sg13g2_decap_8
XFILLER_94_566 VPWR VGND sg13g2_fill_1
XFILLER_48_950 VPWR VGND sg13g2_decap_8
XFILLER_81_238 VPWR VGND sg13g2_decap_8
XFILLER_75_780 VPWR VGND sg13g2_fill_1
XFILLER_74_290 VPWR VGND sg13g2_decap_8
XFILLER_62_430 VPWR VGND sg13g2_decap_8
XFILLER_19_195 VPWR VGND sg13g2_decap_8
X_13929_ VPWR _00480_ net7 VGND sg13g2_inv_1
X_07450_ acc_sub.op_sign_logic0.s_a acc_sub.exp_mant_logic0.a\[15\] net1796 _01442_
+ VPWR VGND sg13g2_mux2_1
XFILLER_62_485 VPWR VGND sg13g2_fill_1
XFILLER_62_474 VPWR VGND sg13g2_decap_8
XFILLER_35_699 VPWR VGND sg13g2_decap_4
XFILLER_34_165 VPWR VGND sg13g2_fill_2
XFILLER_34_154 VPWR VGND sg13g2_decap_8
X_07381_ VPWR _01729_ acc_sub.exp_mant_logic0.a\[12\] VGND sg13g2_inv_1
X_09120_ net1787 _03298_ _03296_ _03301_ VPWR VGND _03300_ sg13g2_nand4_1
XFILLER_89_0 VPWR VGND sg13g2_decap_8
X_09051_ _03237_ _03234_ _03236_ VPWR VGND sg13g2_nand2_1
XFILLER_117_900 VPWR VGND sg13g2_decap_8
X_08002_ fp16_sum_pipe.exp_mant_logic0.a\[2\] _02269_ VPWR VGND sg13g2_inv_4
XFILLER_116_410 VPWR VGND sg13g2_decap_8
XFILLER_117_977 VPWR VGND sg13g2_decap_8
XFILLER_104_605 VPWR VGND sg13g2_decap_4
XFILLER_104_638 VPWR VGND sg13g2_decap_8
XFILLER_103_115 VPWR VGND sg13g2_fill_2
XFILLER_89_316 VPWR VGND sg13g2_decap_8
XFILLER_106_36 VPWR VGND sg13g2_decap_8
XFILLER_106_14 VPWR VGND sg13g2_decap_4
XFILLER_89_349 VPWR VGND sg13g2_fill_2
XFILLER_44_1012 VPWR VGND sg13g2_fill_2
XFILLER_44_1001 VPWR VGND sg13g2_decap_8
X_09953_ _04048_ VPWR _04049_ VGND fp16_res_pipe.exp_mant_logic0.b\[13\] _04047_ sg13g2_o21ai_1
X_08904_ VPWR _03091_ _03089_ VGND sg13g2_inv_1
XFILLER_97_360 VPWR VGND sg13g2_decap_8
XFILLER_85_500 VPWR VGND sg13g2_fill_2
XFILLER_58_725 VPWR VGND sg13g2_decap_8
X_09884_ _01224_ net1767 fp16_res_pipe.reg_add_sub.q\[0\] VPWR VGND sg13g2_nand2b_1
X_08835_ _03022_ _03002_ net1789 VPWR VGND sg13g2_nand2_1
XFILLER_100_844 VPWR VGND sg13g2_decap_8
X_08766_ _02957_ acc_sum.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_inv_2
XFILLER_58_769 VPWR VGND sg13g2_decap_8
XFILLER_122_35 VPWR VGND sg13g2_decap_8
X_07717_ _02024_ net1650 VPWR VGND sg13g2_inv_2
XFILLER_85_588 VPWR VGND sg13g2_decap_8
X_08697_ _02911_ _02756_ _02910_ VPWR VGND sg13g2_xnor2_1
XFILLER_54_975 VPWR VGND sg13g2_fill_2
XFILLER_25_110 VPWR VGND sg13g2_decap_8
XFILLER_53_463 VPWR VGND sg13g2_fill_1
X_07579_ _01892_ VPWR _01893_ VGND _01871_ _01879_ sg13g2_o21ai_1
XFILLER_80_271 VPWR VGND sg13g2_decap_8
XFILLER_13_327 VPWR VGND sg13g2_fill_1
XFILLER_13_349 VPWR VGND sg13g2_decap_8
XFILLER_40_168 VPWR VGND sg13g2_decap_8
X_09318_ _03471_ _03470_ _03389_ VPWR VGND sg13g2_nand2_1
XFILLER_9_309 VPWR VGND sg13g2_fill_2
X_10590_ _04608_ acc_sub.x2\[4\] net1927 VPWR VGND sg13g2_nand2_1
XFILLER_127_708 VPWR VGND sg13g2_decap_8
X_09249_ VPWR _03403_ fp16_res_pipe.op_sign_logic0.mantisa_b\[2\] VGND sg13g2_inv_1
XFILLER_31_21 VPWR VGND sg13g2_decap_8
XFILLER_108_944 VPWR VGND sg13g2_decap_8
X_12260_ _06106_ _06104_ _06105_ VPWR VGND sg13g2_nand2_1
XFILLER_107_454 VPWR VGND sg13g2_fill_2
X_11211_ _02957_ _05176_ _05177_ VPWR VGND sg13g2_nor2_1
X_12191_ _06037_ _06028_ _06036_ VPWR VGND sg13g2_nand2_1
XFILLER_123_925 VPWR VGND sg13g2_decap_8
XFILLER_122_402 VPWR VGND sg13g2_decap_8
X_11142_ _05112_ _05111_ VPWR VGND sg13g2_inv_2
XFILLER_95_319 VPWR VGND sg13g2_fill_2
XFILLER_89_872 VPWR VGND sg13g2_decap_8
X_11073_ _05049_ _05050_ VPWR VGND sg13g2_inv_4
XFILLER_49_725 VPWR VGND sg13g2_decap_8
XFILLER_0_253 VPWR VGND sg13g2_decap_8
XFILLER_1_765 VPWR VGND sg13g2_decap_4
X_14901_ _00702_ VGND VPWR _01421_ acc_sub.op_sign_logic0.mantisa_a\[0\] clknet_leaf_61_clk
+ sg13g2_dfrbpq_1
XFILLER_49_758 VPWR VGND sg13g2_decap_8
X_10024_ _04112_ net1689 _04081_ VPWR VGND sg13g2_nand2_1
X_14832_ _00633_ VGND VPWR _01356_ fpdiv.divider0.remainder_reg\[11\] clknet_leaf_73_clk
+ sg13g2_dfrbpq_1
XFILLER_91_503 VPWR VGND sg13g2_fill_2
XFILLER_76_566 VPWR VGND sg13g2_decap_4
XFILLER_64_706 VPWR VGND sg13g2_decap_8
XFILLER_36_408 VPWR VGND sg13g2_decap_8
XFILLER_64_739 VPWR VGND sg13g2_fill_2
XFILLER_56_62 VPWR VGND sg13g2_decap_8
XFILLER_91_558 VPWR VGND sg13g2_fill_2
X_14763_ _00564_ VGND VPWR _01287_ acc_sum.exp_mant_logic0.b\[8\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
XFILLER_56_290 VPWR VGND sg13g2_fill_1
X_11975_ fpmul.reg_b_out\[11\] fpmul.reg_a_out\[11\] _05829_ VPWR VGND sg13g2_xor2_1
XFILLER_44_441 VPWR VGND sg13g2_decap_8
X_13714_ VPWR _00265_ net58 VGND sg13g2_inv_1
XFILLER_45_997 VPWR VGND sg13g2_decap_4
XFILLER_44_452 VPWR VGND sg13g2_fill_2
X_14694_ _00495_ VGND VPWR _01222_ fp16_res_pipe.op_sign_logic0.s_b clknet_leaf_130_clk
+ sg13g2_dfrbpq_2
XFILLER_16_165 VPWR VGND sg13g2_fill_2
X_10926_ _04849_ _04826_ _04934_ VPWR VGND sg13g2_nor2_1
X_13645_ VPWR _00196_ net111 VGND sg13g2_inv_1
XFILLER_60_967 VPWR VGND sg13g2_fill_2
XFILLER_16_176 VPWR VGND sg13g2_fill_1
X_10857_ VGND VPWR _04806_ net1824 _04869_ _04868_ sg13g2_a21oi_1
XFILLER_72_94 VPWR VGND sg13g2_decap_8
X_13576_ VPWR _00127_ net22 VGND sg13g2_inv_1
XFILLER_9_843 VPWR VGND sg13g2_decap_8
XFILLER_12_360 VPWR VGND sg13g2_decap_8
X_10788_ VPWR _04800_ _04799_ VGND sg13g2_inv_1
XFILLER_31_179 VPWR VGND sg13g2_decap_8
XFILLER_118_719 VPWR VGND sg13g2_decap_8
X_12527_ _06349_ VPWR _00946_ VGND net1956 _05783_ sg13g2_o21ai_1
X_12458_ VPWR _06301_ fpmul.seg_reg0.q\[12\] VGND sg13g2_inv_1
X_11409_ VPWR _05350_ fpdiv.div_out\[2\] VGND sg13g2_inv_1
XFILLER_67_1012 VPWR VGND sg13g2_fill_2
XFILLER_126_785 VPWR VGND sg13g2_decap_8
XFILLER_125_273 VPWR VGND sg13g2_decap_8
XFILLER_99_636 VPWR VGND sg13g2_decap_4
X_12389_ VPWR _06235_ _06229_ VGND sg13g2_inv_1
XFILLER_114_958 VPWR VGND sg13g2_decap_8
XFILLER_98_135 VPWR VGND sg13g2_decap_8
X_14128_ VPWR _00679_ net119 VGND sg13g2_inv_1
XFILLER_4_581 VPWR VGND sg13g2_decap_4
XFILLER_122_980 VPWR VGND sg13g2_decap_8
XFILLER_100_107 VPWR VGND sg13g2_decap_4
XFILLER_97_80 VPWR VGND sg13g2_fill_1
X_14059_ VPWR _00610_ net79 VGND sg13g2_inv_1
XFILLER_100_129 VPWR VGND sg13g2_decap_8
XFILLER_79_382 VPWR VGND sg13g2_fill_1
X_08620_ VPWR _02842_ _02762_ VGND sg13g2_inv_1
XFILLER_55_717 VPWR VGND sg13g2_decap_4
XFILLER_95_897 VPWR VGND sg13g2_fill_1
XFILLER_94_396 VPWR VGND sg13g2_decap_8
XFILLER_94_374 VPWR VGND sg13g2_fill_1
XFILLER_94_363 VPWR VGND sg13g2_decap_8
XFILLER_36_920 VPWR VGND sg13g2_decap_8
X_08551_ VPWR _02775_ _02774_ VGND sg13g2_inv_1
X_07502_ VPWR _01824_ acc_sub.seg_reg0.q\[28\] VGND sg13g2_inv_1
X_08482_ VPWR _02711_ _02710_ VGND sg13g2_inv_1
XFILLER_63_772 VPWR VGND sg13g2_decap_4
XFILLER_36_997 VPWR VGND sg13g2_decap_8
X_07433_ VGND VPWR _01763_ net1749 _01449_ _01765_ sg13g2_a21oi_1
XFILLER_22_124 VPWR VGND sg13g2_fill_2
XFILLER_23_636 VPWR VGND sg13g2_fill_1
XFILLER_23_647 VPWR VGND sg13g2_fill_2
XFILLER_10_308 VPWR VGND sg13g2_decap_8
X_09103_ _03089_ VPWR _03285_ VGND _03180_ _03284_ sg13g2_o21ai_1
X_07364_ _01718_ VPWR _01471_ VGND net1798 _01717_ sg13g2_o21ai_1
XFILLER_10_319 VPWR VGND sg13g2_fill_1
X_07295_ _01662_ _01521_ _01609_ VPWR VGND sg13g2_xnor2_1
XFILLER_108_207 VPWR VGND sg13g2_decap_8
XFILLER_31_691 VPWR VGND sg13g2_decap_8
X_09034_ VPWR _03220_ _03219_ VGND sg13g2_inv_1
XFILLER_117_774 VPWR VGND sg13g2_decap_8
XFILLER_117_35 VPWR VGND sg13g2_decap_8
XFILLER_2_507 VPWR VGND sg13g2_decap_8
XFILLER_105_958 VPWR VGND sg13g2_decap_8
XFILLER_120_939 VPWR VGND sg13g2_decap_8
XFILLER_104_457 VPWR VGND sg13g2_decap_4
X_09936_ VPWR _04032_ fp16_res_pipe.seg_reg0.q\[28\] VGND sg13g2_inv_1
XFILLER_113_991 VPWR VGND sg13g2_decap_8
X_09867_ VGND VPWR _03722_ net1820 _01230_ _03973_ sg13g2_a21oi_1
XFILLER_97_190 VPWR VGND sg13g2_decap_8
XFILLER_86_853 VPWR VGND sg13g2_decap_4
X_09798_ _03663_ VPWR _03912_ VGND _03882_ _03911_ sg13g2_o21ai_1
XFILLER_85_363 VPWR VGND sg13g2_fill_1
Xclkbuf_5_23__f_clk clknet_4_11_0_clk clknet_5_23__leaf_clk VPWR VGND sg13g2_buf_8
X_08749_ _02946_ acc\[9\] net1897 VPWR VGND sg13g2_nand2_1
XFILLER_73_558 VPWR VGND sg13g2_fill_1
XFILLER_73_547 VPWR VGND sg13g2_decap_8
XFILLER_26_21 VPWR VGND sg13g2_decap_8
XFILLER_27_953 VPWR VGND sg13g2_decap_8
X_11760_ _05664_ net1838 fp16_sum_pipe.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_81_580 VPWR VGND sg13g2_decap_8
X_10711_ _04672_ _04723_ _04722_ _04724_ VPWR VGND sg13g2_nand3_1
XFILLER_42_978 VPWR VGND sg13g2_fill_2
XFILLER_41_455 VPWR VGND sg13g2_decap_4
XFILLER_13_146 VPWR VGND sg13g2_decap_4
X_11691_ _05595_ _05583_ _05594_ VPWR VGND sg13g2_nand2_1
X_13430_ _07094_ _07076_ instr\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_42_42 VPWR VGND sg13g2_decap_8
X_10642_ VPWR _04655_ _04652_ VGND sg13g2_inv_1
X_13361_ _07054_ VPWR _00818_ VGND _06941_ _07027_ sg13g2_o21ai_1
X_10573_ _04599_ VPWR _01150_ VGND net1931 _02186_ sg13g2_o21ai_1
XFILLER_10_842 VPWR VGND sg13g2_decap_8
XFILLER_22_691 VPWR VGND sg13g2_fill_2
XFILLER_127_527 VPWR VGND sg13g2_decap_8
X_13292_ _07006_ sipo.word\[4\] VPWR VGND sg13g2_inv_2
X_12312_ _06158_ _05954_ _06067_ VPWR VGND sg13g2_xnor2_1
XFILLER_108_752 VPWR VGND sg13g2_decap_8
X_12243_ _06089_ net1855 net1867 VPWR VGND sg13g2_nand2_1
XFILLER_6_857 VPWR VGND sg13g2_decap_8
XFILLER_123_700 VPWR VGND sg13g2_decap_4
XFILLER_107_251 VPWR VGND sg13g2_decap_8
XFILLER_5_378 VPWR VGND sg13g2_fill_2
XFILLER_122_210 VPWR VGND sg13g2_decap_8
X_12174_ _06018_ _06019_ _05978_ _06020_ VPWR VGND sg13g2_nand3_1
XFILLER_123_799 VPWR VGND sg13g2_decap_8
X_11125_ _05095_ _05094_ _04998_ VPWR VGND sg13g2_nand2_1
XFILLER_3_14 VPWR VGND sg13g2_decap_8
XFILLER_122_287 VPWR VGND sg13g2_decap_4
XFILLER_110_449 VPWR VGND sg13g2_decap_8
X_11056_ _05033_ VPWR _05034_ VGND _05013_ _05032_ sg13g2_o21ai_1
XFILLER_103_490 VPWR VGND sg13g2_decap_4
XFILLER_92_801 VPWR VGND sg13g2_fill_1
XFILLER_88_190 VPWR VGND sg13g2_decap_8
XFILLER_77_853 VPWR VGND sg13g2_decap_4
XFILLER_76_330 VPWR VGND sg13g2_fill_2
X_10007_ _04050_ VPWR _04095_ VGND _04001_ _04094_ sg13g2_o21ai_1
XFILLER_97_1005 VPWR VGND sg13g2_decap_8
XFILLER_18_920 VPWR VGND sg13g2_decap_8
X_14815_ _00616_ VGND VPWR _01339_ acc_sum.add_renorm0.mantisa\[4\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_91_333 VPWR VGND sg13g2_decap_8
XFILLER_45_783 VPWR VGND sg13g2_decap_8
X_14746_ _00547_ VGND VPWR _01274_ fp16_res_pipe.add_renorm0.mantisa\[9\] clknet_leaf_139_clk
+ sg13g2_dfrbpq_2
XFILLER_18_997 VPWR VGND sg13g2_decap_8
XFILLER_91_399 VPWR VGND sg13g2_decap_8
X_11958_ _05816_ net1883 fpmul.reg_b_out\[3\] VPWR VGND sg13g2_nand2_1
X_11889_ _05775_ VPWR _01010_ VGND _05774_ _05767_ sg13g2_o21ai_1
XFILLER_60_775 VPWR VGND sg13g2_decap_8
XFILLER_44_293 VPWR VGND sg13g2_decap_8
XFILLER_33_967 VPWR VGND sg13g2_decap_8
X_14677_ _00478_ VGND VPWR _01205_ fp16_res_pipe.op_sign_logic0.mantisa_a\[3\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_10909_ _04737_ VPWR _04918_ VGND _04903_ _04917_ sg13g2_o21ai_1
X_13628_ VPWR _00179_ net57 VGND sg13g2_inv_1
X_13559_ VPWR _00110_ net21 VGND sg13g2_inv_1
XFILLER_8_161 VPWR VGND sg13g2_decap_8
XFILLER_114_755 VPWR VGND sg13g2_decap_8
XFILLER_99_444 VPWR VGND sg13g2_decap_8
Xfanout107 net141 net107 VPWR VGND sg13g2_buf_2
Xfanout129 net140 net129 VPWR VGND sg13g2_buf_2
XFILLER_87_628 VPWR VGND sg13g2_decap_8
Xfanout118 net119 net118 VPWR VGND sg13g2_buf_2
X_07982_ _02254_ fp16_sum_pipe.exp_mant_logic0.a\[11\] _02250_ fp16_sum_pipe.seg_reg0.q\[26\]
+ net1775 VPWR VGND sg13g2_a22oi_1
XFILLER_113_287 VPWR VGND sg13g2_decap_4
X_09721_ _03834_ _03836_ _03837_ VPWR VGND sg13g2_nor2_1
XFILLER_101_416 VPWR VGND sg13g2_decap_8
XFILLER_99_499 VPWR VGND sg13g2_fill_1
XFILLER_68_864 VPWR VGND sg13g2_fill_1
XFILLER_110_983 VPWR VGND sg13g2_decap_8
X_09652_ _03769_ _03674_ _03661_ _03649_ _03635_ VPWR VGND sg13g2_a22oi_1
XFILLER_55_514 VPWR VGND sg13g2_fill_1
X_09583_ VGND VPWR _02806_ acc_sum.add_renorm0.mantisa\[4\] _03700_ _03699_ sg13g2_a21oi_1
XFILLER_83_845 VPWR VGND sg13g2_decap_8
X_08603_ VGND VPWR _02823_ _02758_ _02826_ _02825_ sg13g2_a21oi_1
XFILLER_55_547 VPWR VGND sg13g2_fill_1
XFILLER_27_227 VPWR VGND sg13g2_decap_4
X_08534_ VPWR _02758_ _02753_ VGND sg13g2_inv_1
XFILLER_42_219 VPWR VGND sg13g2_decap_8
XFILLER_35_260 VPWR VGND sg13g2_decap_8
X_08465_ _01356_ net1718 _02697_ _02652_ _02689_ VPWR VGND sg13g2_a22oi_1
XFILLER_51_742 VPWR VGND sg13g2_decap_8
XFILLER_24_967 VPWR VGND sg13g2_decap_8
X_07416_ _01752_ VPWR _01453_ VGND net1894 _01751_ sg13g2_o21ai_1
X_08396_ _02633_ _02618_ _02569_ VPWR VGND sg13g2_nand2_1
XFILLER_10_105 VPWR VGND sg13g2_decap_8
X_07347_ VPWR _01707_ acc_sub.add_renorm0.mantisa\[0\] VGND sg13g2_inv_1
X_09017_ _03173_ _03094_ _03203_ VPWR VGND sg13g2_xor2_1
X_07278_ _01640_ _01646_ _01639_ _01485_ VPWR VGND sg13g2_nand3_1
XFILLER_12_56 VPWR VGND sg13g2_decap_8
XFILLER_117_560 VPWR VGND sg13g2_fill_1
XFILLER_2_304 VPWR VGND sg13g2_fill_1
XFILLER_117_593 VPWR VGND sg13g2_fill_2
XFILLER_78_606 VPWR VGND sg13g2_decap_4
XFILLER_120_736 VPWR VGND sg13g2_decap_8
XFILLER_120_725 VPWR VGND sg13g2_fill_1
XFILLER_104_287 VPWR VGND sg13g2_fill_2
XFILLER_77_116 VPWR VGND sg13g2_fill_1
XFILLER_59_853 VPWR VGND sg13g2_fill_1
X_09919_ _04013_ _04015_ _04016_ VPWR VGND sg13g2_nor2_1
XFILLER_101_983 VPWR VGND sg13g2_decap_8
XFILLER_86_694 VPWR VGND sg13g2_fill_2
X_12930_ _06702_ _06703_ _06693_ _00898_ VPWR VGND sg13g2_nand3_1
XFILLER_74_834 VPWR VGND sg13g2_decap_8
XFILLER_58_352 VPWR VGND sg13g2_fill_2
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_73_344 VPWR VGND sg13g2_fill_1
X_12861_ VGND VPWR acc\[9\] net1907 _06640_ net1909 sg13g2_a21oi_1
XFILLER_46_569 VPWR VGND sg13g2_fill_2
X_14600_ _00401_ VGND VPWR _01132_ fp16_res_pipe.y\[11\] clknet_leaf_129_clk sg13g2_dfrbpq_2
X_11812_ _05713_ _05712_ _05622_ VPWR VGND sg13g2_nand2_1
X_12792_ _06577_ net1716 _00020_ VPWR VGND sg13g2_nand2_1
XFILLER_14_411 VPWR VGND sg13g2_fill_1
XFILLER_15_945 VPWR VGND sg13g2_decap_8
X_14531_ _00332_ VGND VPWR _01067_ fpdiv.div_out\[6\] clknet_leaf_77_clk sg13g2_dfrbpq_2
XFILLER_42_764 VPWR VGND sg13g2_fill_2
X_11743_ _05587_ _05628_ _05642_ _05647_ VPWR VGND _05610_ sg13g2_nand4_1
XFILLER_14_444 VPWR VGND sg13g2_decap_8
XFILLER_26_293 VPWR VGND sg13g2_decap_8
X_14462_ _00263_ VGND VPWR _01001_ fpmul.seg_reg0.q\[47\] clknet_leaf_125_clk sg13g2_dfrbpq_1
X_11674_ _05578_ _05577_ fp16_sum_pipe.add_renorm0.exp\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_30_948 VPWR VGND sg13g2_decap_8
X_13413_ _07085_ VPWR _00797_ VGND _07037_ net1722 sg13g2_o21ai_1
X_10625_ _04627_ _04637_ _04638_ VPWR VGND sg13g2_nor2_1
X_14393_ _00194_ VGND VPWR _00932_ div_result\[6\] clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_127_357 VPWR VGND sg13g2_decap_8
X_13344_ _07045_ VPWR _00826_ VGND _07044_ net1726 sg13g2_o21ai_1
X_10556_ _04589_ fp16_sum_pipe.add_renorm0.exp\[3\] VPWR VGND sg13g2_inv_2
X_13275_ _06993_ net1729 acc_sum.y\[8\] VPWR VGND sg13g2_nand2_1
X_10487_ _04493_ VPWR _04533_ VGND _04531_ _04532_ sg13g2_o21ai_1
XFILLER_108_582 VPWR VGND sg13g2_decap_8
X_12226_ _06072_ net1855 net1868 VPWR VGND sg13g2_nand2_1
XFILLER_45_7 VPWR VGND sg13g2_decap_8
XFILLER_5_175 VPWR VGND sg13g2_decap_4
XFILLER_69_606 VPWR VGND sg13g2_fill_2
X_12157_ _06003_ _06002_ _05987_ VPWR VGND sg13g2_nand2b_1
XFILLER_123_574 VPWR VGND sg13g2_decap_8
XFILLER_111_747 VPWR VGND sg13g2_decap_8
XFILLER_111_736 VPWR VGND sg13g2_fill_1
XFILLER_110_213 VPWR VGND sg13g2_fill_1
XFILLER_96_425 VPWR VGND sg13g2_decap_8
X_11108_ _05077_ VPWR _05078_ VGND _05022_ _05019_ sg13g2_o21ai_1
XFILLER_77_650 VPWR VGND sg13g2_decap_8
X_12088_ _05899_ _05900_ _05934_ VPWR VGND sg13g2_nor2_1
XFILLER_49_330 VPWR VGND sg13g2_decap_8
X_11039_ _05018_ _05014_ _05017_ VPWR VGND sg13g2_nand2_1
XFILLER_49_363 VPWR VGND sg13g2_decap_8
XFILLER_92_620 VPWR VGND sg13g2_fill_1
XFILLER_49_396 VPWR VGND sg13g2_decap_8
XFILLER_92_675 VPWR VGND sg13g2_fill_1
XFILLER_80_826 VPWR VGND sg13g2_decap_4
XFILLER_65_889 VPWR VGND sg13g2_decap_8
XFILLER_64_377 VPWR VGND sg13g2_fill_2
XFILLER_24_208 VPWR VGND sg13g2_fill_1
XFILLER_64_388 VPWR VGND sg13g2_decap_4
XFILLER_45_591 VPWR VGND sg13g2_decap_8
XFILLER_45_580 VPWR VGND sg13g2_decap_8
X_14729_ _00530_ VGND VPWR _01257_ fp16_res_pipe.add_renorm0.exp\[0\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_2
XFILLER_60_583 VPWR VGND sg13g2_decap_8
X_08250_ _02501_ fp16_sum_pipe.exp_mant_logic0.b\[3\] net1645 _02472_ net1657 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_32_274 VPWR VGND sg13g2_decap_8
X_07201_ VGND VPWR _01572_ _01538_ _01573_ _01532_ sg13g2_a21oi_1
XFILLER_119_814 VPWR VGND sg13g2_decap_8
X_08181_ _02261_ _02427_ _02439_ VPWR VGND sg13g2_nor2_1
XFILLER_20_447 VPWR VGND sg13g2_decap_8
XFILLER_21_959 VPWR VGND sg13g2_decap_8
X_07132_ acc_sub.op_sign_logic0.mantisa_b\[8\] _01503_ _01504_ VPWR VGND sg13g2_nor2_1
XFILLER_71_0 VPWR VGND sg13g2_decap_4
XFILLER_106_519 VPWR VGND sg13g2_decap_8
XFILLER_114_530 VPWR VGND sg13g2_decap_8
XFILLER_99_241 VPWR VGND sg13g2_decap_8
XFILLER_99_296 VPWR VGND sg13g2_decap_8
XFILLER_114_14 VPWR VGND sg13g2_decap_8
X_07965_ fp16_sum_pipe.exp_mant_logic0.b\[14\] _02238_ _02239_ VPWR VGND sg13g2_nor2_1
X_09704_ _03820_ acc_sum.add_renorm0.exp\[6\] _03791_ VPWR VGND sg13g2_xnor2_1
XFILLER_68_683 VPWR VGND sg13g2_decap_8
XFILLER_110_780 VPWR VGND sg13g2_decap_8
X_09635_ _03752_ _03649_ _03655_ VPWR VGND sg13g2_nand2_1
X_07896_ _02175_ net1891 acc_sub.x2\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_56_856 VPWR VGND sg13g2_decap_8
XFILLER_55_355 VPWR VGND sg13g2_decap_4
X_09566_ net1803 VPWR _03683_ VGND _03665_ _03681_ sg13g2_o21ai_1
XFILLER_82_174 VPWR VGND sg13g2_fill_2
XFILLER_43_539 VPWR VGND sg13g2_decap_8
XFILLER_36_580 VPWR VGND sg13g2_decap_8
X_08517_ _02741_ _02739_ acc_sum.op_sign_logic0.mantisa_b\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_70_347 VPWR VGND sg13g2_fill_2
XFILLER_12_904 VPWR VGND sg13g2_decap_8
XFILLER_23_230 VPWR VGND sg13g2_decap_4
XFILLER_24_764 VPWR VGND sg13g2_fill_2
X_09497_ _03616_ acc_sub.x2\[1\] net1916 VPWR VGND sg13g2_nand2_1
X_08448_ _02682_ _02679_ fpdiv.divider0.divisor_reg\[11\] _02680_ VPWR VGND sg13g2_and3_1
XFILLER_51_572 VPWR VGND sg13g2_decap_8
XFILLER_23_274 VPWR VGND sg13g2_fill_2
X_08379_ _02620_ _07115_ fpdiv.reg2en.q\[0\] VPWR VGND sg13g2_nand2b_1
XFILLER_7_418 VPWR VGND sg13g2_fill_2
XFILLER_7_407 VPWR VGND sg13g2_fill_1
X_10410_ VGND VPWR _04459_ _04460_ _04458_ _04456_ sg13g2_a21oi_2
XFILLER_23_77 VPWR VGND sg13g2_decap_8
XFILLER_99_15 VPWR VGND sg13g2_fill_1
X_11390_ _05338_ VPWR _01072_ VGND _05337_ net1706 sg13g2_o21ai_1
X_10341_ _04391_ _04390_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_118_880 VPWR VGND sg13g2_decap_8
X_13060_ VPWR _06828_ _06827_ VGND sg13g2_inv_1
XFILLER_3_646 VPWR VGND sg13g2_decap_8
XFILLER_2_112 VPWR VGND sg13g2_decap_8
X_10272_ _04341_ VPWR _04342_ VGND _04298_ _04233_ sg13g2_o21ai_1
XFILLER_117_390 VPWR VGND sg13g2_fill_1
XFILLER_79_915 VPWR VGND sg13g2_decap_8
X_12011_ _05863_ fpmul.seg_reg0.q\[21\] VPWR VGND sg13g2_inv_2
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_94_907 VPWR VGND sg13g2_fill_2
XFILLER_120_588 VPWR VGND sg13g2_fill_2
XFILLER_120_566 VPWR VGND sg13g2_decap_4
XFILLER_93_428 VPWR VGND sg13g2_decap_8
X_13962_ VPWR _00513_ net79 VGND sg13g2_inv_1
XFILLER_59_683 VPWR VGND sg13g2_decap_8
XFILLER_58_160 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_111_1013 VPWR VGND sg13g2_fill_1
X_12913_ VPWR _06688_ fpmul.reg_p_out\[5\] VGND sg13g2_inv_1
XFILLER_46_333 VPWR VGND sg13g2_decap_8
XFILLER_74_675 VPWR VGND sg13g2_decap_8
XFILLER_73_130 VPWR VGND sg13g2_decap_4
X_13893_ VPWR _00444_ net35 VGND sg13g2_inv_1
X_12844_ _06625_ net1716 _00016_ VPWR VGND sg13g2_nand2_1
XFILLER_61_303 VPWR VGND sg13g2_fill_1
XFILLER_46_388 VPWR VGND sg13g2_fill_2
XFILLER_64_95 VPWR VGND sg13g2_decap_4
XFILLER_61_369 VPWR VGND sg13g2_decap_4
X_14514_ _00315_ VGND VPWR _01050_ fpdiv.divider0.dividend\[9\] clknet_leaf_58_clk
+ sg13g2_dfrbpq_1
X_11726_ _05630_ _05587_ _05629_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_35 VPWR VGND sg13g2_decap_8
XFILLER_15_797 VPWR VGND sg13g2_fill_2
XFILLER_80_50 VPWR VGND sg13g2_decap_8
X_14445_ _00246_ VGND VPWR _00984_ fpmul.seg_reg0.q\[30\] clknet_leaf_103_clk sg13g2_dfrbpq_1
X_11657_ VGND VPWR _05559_ net1837 _05562_ _05561_ sg13g2_a21oi_1
X_14376_ _00177_ VGND VPWR _00917_ fpmul.reg_b_out\[7\] clknet_leaf_96_clk sg13g2_dfrbpq_2
XFILLER_7_930 VPWR VGND sg13g2_decap_8
X_10608_ _04621_ fp16_res_pipe.add_renorm0.mantisa\[5\] VPWR VGND sg13g2_inv_2
X_11588_ _05493_ _05457_ _05492_ VPWR VGND sg13g2_nand2_2
XFILLER_127_154 VPWR VGND sg13g2_decap_8
XFILLER_116_828 VPWR VGND sg13g2_decap_8
X_13327_ VPWR _07034_ sipo.word\[13\] VGND sg13g2_inv_1
X_10539_ net1849 fp16_sum_pipe.add_renorm0.mantisa\[1\] _04578_ VPWR VGND sg13g2_nor2_1
XFILLER_115_327 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_decap_8
XFILLER_124_872 VPWR VGND sg13g2_decap_8
X_13258_ _06980_ sipo.word\[12\] VPWR VGND sg13g2_inv_2
XFILLER_9_1004 VPWR VGND sg13g2_decap_8
X_12209_ VGND VPWR _06013_ _06016_ _06055_ _06054_ sg13g2_a21oi_1
X_13189_ VPWR _06927_ sipo.shift_reg\[8\] VGND sg13g2_inv_1
X_07750_ acc_sub.exp_mant_logic0.b\[10\] acc_sub.exp_mant_logic0.b\[9\] acc_sub.exp_mant_logic0.b\[8\]
+ acc_sub.exp_mant_logic0.b\[7\] _02054_ VPWR VGND sg13g2_nor4_1
XFILLER_85_929 VPWR VGND sg13g2_decap_8
XFILLER_78_992 VPWR VGND sg13g2_decap_4
XFILLER_78_981 VPWR VGND sg13g2_decap_4
XFILLER_38_823 VPWR VGND sg13g2_fill_2
XFILLER_93_940 VPWR VGND sg13g2_decap_8
XFILLER_38_834 VPWR VGND sg13g2_decap_8
XFILLER_80_612 VPWR VGND sg13g2_fill_1
X_09420_ _03564_ _03562_ _03563_ fp16_res_pipe.add_renorm0.mantisa\[2\] net1770 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_18_580 VPWR VGND sg13g2_decap_4
X_09351_ _03485_ _03502_ _03484_ _01275_ VPWR VGND sg13g2_nand3_1
X_09282_ _03371_ _03435_ _03436_ VPWR VGND sg13g2_nor2_2
X_08302_ _02545_ _02548_ _02544_ _02549_ VPWR VGND sg13g2_nand3_1
XFILLER_33_550 VPWR VGND sg13g2_decap_8
XFILLER_61_892 VPWR VGND sg13g2_fill_2
X_08233_ _02486_ net1645 net1842 VPWR VGND sg13g2_nand2_1
XFILLER_20_233 VPWR VGND sg13g2_fill_1
XFILLER_109_14 VPWR VGND sg13g2_decap_8
X_08164_ _02422_ VPWR _02423_ VGND _02269_ net1648 sg13g2_o21ai_1
XFILLER_118_154 VPWR VGND sg13g2_decap_8
X_08095_ _02358_ _02359_ _02356_ _02360_ VPWR VGND sg13g2_nand3_1
Xclkload70 VPWR clkload70/Y clknet_leaf_30_clk VGND sg13g2_inv_1
Xclkload81 clkload81/Y clknet_leaf_38_clk VPWR VGND sg13g2_inv_2
XFILLER_88_701 VPWR VGND sg13g2_fill_2
Xclkload92 clkload92/Y clknet_leaf_89_clk VPWR VGND sg13g2_inv_2
XFILLER_115_872 VPWR VGND sg13g2_decap_8
XFILLER_88_734 VPWR VGND sg13g2_fill_1
XFILLER_88_723 VPWR VGND sg13g2_decap_8
XFILLER_125_35 VPWR VGND sg13g2_decap_8
XFILLER_87_244 VPWR VGND sg13g2_fill_2
X_08997_ VGND VPWR _03182_ _03183_ _03145_ _01713_ sg13g2_a21oi_2
XFILLER_88_789 VPWR VGND sg13g2_decap_8
XFILLER_87_277 VPWR VGND sg13g2_decap_8
XFILLER_69_970 VPWR VGND sg13g2_decap_8
XFILLER_29_801 VPWR VGND sg13g2_decap_4
XFILLER_102_599 VPWR VGND sg13g2_fill_1
XFILLER_56_620 VPWR VGND sg13g2_decap_8
X_07948_ _02223_ _02202_ _02222_ VPWR VGND sg13g2_nand2_2
XFILLER_84_973 VPWR VGND sg13g2_decap_8
X_07879_ _02166_ VPWR _01404_ VGND net1885 _01804_ sg13g2_o21ai_1
XFILLER_56_675 VPWR VGND sg13g2_decap_4
XFILLER_56_664 VPWR VGND sg13g2_decap_8
XFILLER_28_355 VPWR VGND sg13g2_decap_8
X_09618_ _03735_ _03723_ _03729_ VPWR VGND sg13g2_xnor2_1
XFILLER_71_623 VPWR VGND sg13g2_fill_2
XFILLER_70_111 VPWR VGND sg13g2_decap_8
XFILLER_55_163 VPWR VGND sg13g2_decap_8
X_10890_ _04901_ _04772_ fp16_res_pipe.y\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_16_528 VPWR VGND sg13g2_decap_8
XFILLER_16_539 VPWR VGND sg13g2_fill_1
X_09549_ _03644_ _03630_ _03666_ VPWR VGND sg13g2_nor2_2
XFILLER_34_21 VPWR VGND sg13g2_decap_8
XFILLER_70_155 VPWR VGND sg13g2_fill_2
XFILLER_52_881 VPWR VGND sg13g2_fill_1
X_12560_ _06376_ fpdiv.reg_a_out\[8\] fpdiv.reg_b_out\[8\] VPWR VGND sg13g2_xnor2_1
XFILLER_34_98 VPWR VGND sg13g2_decap_8
X_12491_ _06241_ _06224_ _06327_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_705 VPWR VGND sg13g2_decap_8
XFILLER_11_266 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_decap_8
X_11511_ _05412_ _05415_ _05416_ VPWR VGND sg13g2_nor2_1
X_11442_ _05371_ acc_sub.x2\[7\] fpdiv.reg1en.d\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_50_42 VPWR VGND sg13g2_decap_8
X_14230_ _00031_ VGND VPWR _00781_ sipo.shift_reg\[11\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_7_226 VPWR VGND sg13g2_decap_8
XFILLER_119_0 VPWR VGND sg13g2_decap_8
X_14161_ VPWR _00712_ net132 VGND sg13g2_inv_1
X_11373_ _05321_ _05322_ _05323_ _05324_ VPWR VGND sg13g2_nor3_1
XFILLER_109_187 VPWR VGND sg13g2_fill_2
X_13112_ _06779_ _06868_ _06869_ VPWR VGND sg13g2_nor2_1
XFILLER_4_944 VPWR VGND sg13g2_decap_8
X_10324_ _04379_ VPWR _01179_ VGND net1921 _04300_ sg13g2_o21ai_1
XFILLER_113_809 VPWR VGND sg13g2_decap_8
X_14092_ VPWR _00643_ net40 VGND sg13g2_inv_1
XFILLER_124_168 VPWR VGND sg13g2_decap_8
XFILLER_79_712 VPWR VGND sg13g2_decap_8
X_13043_ VPWR _06811_ _06810_ VGND sg13g2_inv_1
XFILLER_3_476 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
X_10255_ _04326_ _04210_ net1745 VPWR VGND sg13g2_nand2_1
XFILLER_105_393 VPWR VGND sg13g2_decap_4
XFILLER_59_73 VPWR VGND sg13g2_fill_2
X_10186_ fp16_res_pipe.exp_mant_logic0.b\[10\] fp16_res_pipe.exp_mant_logic0.b\[9\]
+ fp16_res_pipe.exp_mant_logic0.b\[8\] fp16_res_pipe.exp_mant_logic0.b\[7\] _04264_
+ VPWR VGND sg13g2_nor4_1
XFILLER_121_875 VPWR VGND sg13g2_decap_8
XFILLER_120_363 VPWR VGND sg13g2_fill_2
XFILLER_38_119 VPWR VGND sg13g2_decap_8
XFILLER_94_759 VPWR VGND sg13g2_decap_8
XFILLER_93_236 VPWR VGND sg13g2_decap_8
XFILLER_59_491 VPWR VGND sg13g2_decap_8
XFILLER_19_300 VPWR VGND sg13g2_decap_8
XFILLER_93_269 VPWR VGND sg13g2_decap_8
XFILLER_75_50 VPWR VGND sg13g2_decap_4
XFILLER_47_675 VPWR VGND sg13g2_decap_8
X_13945_ VPWR _00496_ net27 VGND sg13g2_inv_1
XFILLER_90_932 VPWR VGND sg13g2_decap_8
XFILLER_90_921 VPWR VGND sg13g2_fill_1
XFILLER_75_995 VPWR VGND sg13g2_decap_8
XFILLER_75_94 VPWR VGND sg13g2_decap_8
X_13876_ VPWR _00427_ net53 VGND sg13g2_inv_1
X_12827_ _06609_ _06605_ _06608_ _06485_ net1941 VPWR VGND sg13g2_a22oi_1
XFILLER_43_881 VPWR VGND sg13g2_decap_8
XFILLER_15_572 VPWR VGND sg13g2_decap_8
XFILLER_61_188 VPWR VGND sg13g2_decap_4
X_12758_ _06545_ VPWR _00912_ VGND net1957 _06015_ sg13g2_o21ai_1
XFILLER_43_892 VPWR VGND sg13g2_decap_8
X_12689_ VPWR _06499_ div_result\[8\] VGND sg13g2_inv_1
X_11709_ _05613_ _05612_ _04583_ VPWR VGND sg13g2_nand2_1
X_14428_ _00229_ VGND VPWR _00967_ fpmul.seg_reg0.q\[13\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_7_760 VPWR VGND sg13g2_decap_8
XFILLER_116_636 VPWR VGND sg13g2_fill_2
X_14359_ _00160_ VGND VPWR _00901_ _00012_ clknet_leaf_87_clk sg13g2_dfrbpq_1
Xfanout9 net10 net9 VPWR VGND sg13g2_buf_2
X_08920_ _03107_ _02971_ _03017_ _03014_ _02996_ VPWR VGND sg13g2_a22oi_1
XFILLER_115_168 VPWR VGND sg13g2_decap_8
XFILLER_103_319 VPWR VGND sg13g2_fill_2
XFILLER_97_520 VPWR VGND sg13g2_fill_2
XFILLER_69_211 VPWR VGND sg13g2_decap_8
X_08851_ _03037_ VPWR _03038_ VGND net1789 _02975_ sg13g2_o21ai_1
XFILLER_112_831 VPWR VGND sg13g2_decap_8
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_07802_ _02101_ acc_sub.exp_mant_logic0.b\[2\] net1669 acc_sub.op_sign_logic0.mantisa_b\[5\]
+ net1779 VPWR VGND sg13g2_a22oi_1
XFILLER_85_726 VPWR VGND sg13g2_decap_8
XFILLER_58_918 VPWR VGND sg13g2_decap_8
X_08782_ VPWR _02969_ _02966_ VGND sg13g2_inv_1
XFILLER_111_374 VPWR VGND sg13g2_fill_2
XFILLER_84_236 VPWR VGND sg13g2_fill_1
XFILLER_66_940 VPWR VGND sg13g2_decap_8
XFILLER_38_631 VPWR VGND sg13g2_decap_8
X_07733_ _02037_ _02038_ _02039_ VPWR VGND _02032_ sg13g2_nand3b_1
XFILLER_84_247 VPWR VGND sg13g2_decap_8
Xclkbuf_5_4__f_clk clknet_4_2_0_clk clknet_5_4__leaf_clk VPWR VGND sg13g2_buf_8
X_07664_ _01910_ _01933_ _01974_ VPWR VGND sg13g2_nor2_1
XFILLER_38_697 VPWR VGND sg13g2_decap_8
XFILLER_37_152 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_92_280 VPWR VGND sg13g2_fill_1
XFILLER_37_196 VPWR VGND sg13g2_fill_2
X_09403_ _03546_ _03548_ _03545_ _01269_ VPWR VGND sg13g2_nand3_1
X_07595_ VPWR _01909_ _01908_ VGND sg13g2_inv_1
XFILLER_80_464 VPWR VGND sg13g2_decap_8
XFILLER_80_453 VPWR VGND sg13g2_fill_2
XFILLER_53_678 VPWR VGND sg13g2_decap_8
XFILLER_52_144 VPWR VGND sg13g2_decap_4
X_09334_ _03375_ VPWR _03486_ VGND fp16_res_pipe.op_sign_logic0.mantisa_a\[8\] _03434_
+ sg13g2_o21ai_1
X_09265_ VGND VPWR _03418_ _03406_ _03419_ _03401_ sg13g2_a21oi_1
X_09196_ _03354_ acc_sub.x2\[2\] net1906 VPWR VGND sg13g2_nand2_1
X_08216_ _02471_ _02472_ VPWR VGND sg13g2_inv_4
XFILLER_119_441 VPWR VGND sg13g2_fill_2
XFILLER_112_7 VPWR VGND sg13g2_decap_8
X_08147_ _02341_ _02327_ _02407_ VPWR VGND sg13g2_nor2_1
XFILLER_20_56 VPWR VGND sg13g2_decap_8
XFILLER_121_105 VPWR VGND sg13g2_decap_8
Xplace1960 net1959 net1960 VPWR VGND sg13g2_buf_1
XFILLER_96_49 VPWR VGND sg13g2_fill_2
XFILLER_88_553 VPWR VGND sg13g2_fill_2
XFILLER_88_520 VPWR VGND sg13g2_fill_1
XFILLER_0_435 VPWR VGND sg13g2_decap_8
XFILLER_1_969 VPWR VGND sg13g2_decap_8
X_10040_ _04114_ _04120_ _04128_ VPWR VGND sg13g2_nor2_2
XFILLER_76_726 VPWR VGND sg13g2_fill_2
XFILLER_29_21 VPWR VGND sg13g2_decap_8
XFILLER_48_428 VPWR VGND sg13g2_decap_8
XFILLER_29_620 VPWR VGND sg13g2_decap_8
XFILLER_63_409 VPWR VGND sg13g2_decap_4
X_11991_ VGND VPWR _05839_ _05843_ _05845_ _05844_ sg13g2_a21oi_1
XFILLER_90_228 VPWR VGND sg13g2_fill_1
X_13730_ VPWR _00281_ net64 VGND sg13g2_inv_1
X_10942_ net1771 VPWR _04949_ VGND _04948_ _04871_ sg13g2_o21ai_1
XFILLER_29_686 VPWR VGND sg13g2_decap_8
XFILLER_90_239 VPWR VGND sg13g2_fill_2
XFILLER_45_42 VPWR VGND sg13g2_decap_8
XFILLER_43_133 VPWR VGND sg13g2_decap_8
X_13661_ VPWR _00212_ net57 VGND sg13g2_inv_1
XFILLER_43_155 VPWR VGND sg13g2_decap_8
XFILLER_25_870 VPWR VGND sg13g2_fill_1
XFILLER_31_306 VPWR VGND sg13g2_decap_8
X_10873_ VPWR _04884_ _04813_ VGND sg13g2_inv_1
XFILLER_32_818 VPWR VGND sg13g2_decap_8
XFILLER_101_70 VPWR VGND sg13g2_decap_4
X_12612_ _06423_ _06427_ _06428_ VPWR VGND sg13g2_nor2_1
X_13592_ VPWR _00143_ net121 VGND sg13g2_inv_1
XFILLER_71_497 VPWR VGND sg13g2_decap_8
XFILLER_24_380 VPWR VGND sg13g2_fill_1
X_12543_ fpdiv.divider0.dividend\[5\] _06355_ _06356_ _06360_ VGND VPWR _06359_ sg13g2_nor4_2
XFILLER_8_513 VPWR VGND sg13g2_fill_1
XFILLER_12_542 VPWR VGND sg13g2_decap_4
XFILLER_8_535 VPWR VGND sg13g2_decap_4
X_14213_ VPWR _00764_ net135 VGND sg13g2_inv_1
X_12474_ _06314_ net1871 _06308_ _06315_ VPWR VGND sg13g2_nand3_1
XFILLER_6_14 VPWR VGND sg13g2_decap_8
XFILLER_125_422 VPWR VGND sg13g2_decap_8
XFILLER_125_411 VPWR VGND sg13g2_fill_1
X_11425_ net1940 fpdiv.reg_a_out\[13\] _05360_ VPWR VGND sg13g2_nor2_1
XFILLER_126_967 VPWR VGND sg13g2_decap_8
X_14144_ VPWR _00695_ net129 VGND sg13g2_inv_1
X_11356_ _01076_ _05307_ _05308_ VPWR VGND sg13g2_nand2_1
XFILLER_112_105 VPWR VGND sg13g2_fill_2
X_14075_ VPWR _00626_ net138 VGND sg13g2_inv_1
X_10307_ _04371_ net1914 fp16_res_pipe.x2\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_106_691 VPWR VGND sg13g2_decap_4
X_13026_ VPWR _06794_ _06793_ VGND sg13g2_inv_1
X_11287_ _01084_ _05246_ _05247_ VPWR VGND sg13g2_nand2_1
X_10238_ _04298_ _04124_ _04310_ VPWR VGND sg13g2_nor2_1
XFILLER_120_182 VPWR VGND sg13g2_decap_8
XFILLER_94_534 VPWR VGND sg13g2_decap_4
XFILLER_67_737 VPWR VGND sg13g2_decap_4
X_10169_ _03617_ _04156_ _04249_ VPWR VGND sg13g2_nor2_1
XFILLER_66_258 VPWR VGND sg13g2_fill_2
XFILLER_47_450 VPWR VGND sg13g2_fill_2
XFILLER_19_141 VPWR VGND sg13g2_decap_8
XFILLER_94_589 VPWR VGND sg13g2_fill_1
XFILLER_81_206 VPWR VGND sg13g2_decap_4
X_13928_ VPWR _00479_ net5 VGND sg13g2_inv_1
XFILLER_19_163 VPWR VGND sg13g2_fill_1
XFILLER_90_751 VPWR VGND sg13g2_fill_1
XFILLER_47_494 VPWR VGND sg13g2_decap_8
XFILLER_35_656 VPWR VGND sg13g2_decap_8
XFILLER_34_133 VPWR VGND sg13g2_decap_8
X_13859_ VPWR _00410_ net14 VGND sg13g2_inv_1
XFILLER_23_807 VPWR VGND sg13g2_fill_1
XFILLER_96_2 VPWR VGND sg13g2_fill_1
X_07380_ _01728_ VPWR _01465_ VGND net1887 _01727_ sg13g2_o21ai_1
XFILLER_34_177 VPWR VGND sg13g2_decap_8
XFILLER_22_317 VPWR VGND sg13g2_decap_8
XFILLER_124_1012 VPWR VGND sg13g2_fill_2
XFILLER_31_851 VPWR VGND sg13g2_decap_8
XFILLER_31_873 VPWR VGND sg13g2_decap_8
X_09050_ _03235_ VPWR _03236_ VGND net1791 _01713_ sg13g2_o21ai_1
X_08001_ _02268_ fp16_sum_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_inv_2
XFILLER_116_400 VPWR VGND sg13g2_decap_4
XFILLER_117_956 VPWR VGND sg13g2_decap_8
XFILLER_7_590 VPWR VGND sg13g2_fill_1
X_09952_ VGND VPWR _04047_ _03591_ _04048_ net1766 sg13g2_a21oi_1
XFILLER_98_840 VPWR VGND sg13g2_decap_8
XFILLER_100_812 VPWR VGND sg13g2_decap_8
XFILLER_100_801 VPWR VGND sg13g2_fill_2
X_08834_ _03020_ VPWR _03021_ VGND net1788 _01647_ sg13g2_o21ai_1
XFILLER_111_182 VPWR VGND sg13g2_fill_2
XFILLER_122_14 VPWR VGND sg13g2_decap_8
X_08765_ _02956_ VPWR _01315_ VGND net1899 _02955_ sg13g2_o21ai_1
XFILLER_73_707 VPWR VGND sg13g2_fill_2
X_07716_ _02022_ VPWR _02023_ VGND _01753_ _01979_ sg13g2_o21ai_1
XFILLER_66_792 VPWR VGND sg13g2_fill_1
XFILLER_39_984 VPWR VGND sg13g2_decap_8
XFILLER_26_612 VPWR VGND sg13g2_decap_8
X_08696_ _02910_ _02908_ _02909_ _02907_ net1739 VPWR VGND sg13g2_a22oi_1
XFILLER_82_18 VPWR VGND sg13g2_fill_1
XFILLER_65_280 VPWR VGND sg13g2_fill_2
XFILLER_53_431 VPWR VGND sg13g2_decap_8
X_07647_ _01929_ net1660 _01959_ VPWR VGND sg13g2_nor2_2
XFILLER_81_784 VPWR VGND sg13g2_decap_4
X_07578_ _01892_ net1687 _01891_ VPWR VGND sg13g2_nand2b_1
XFILLER_80_294 VPWR VGND sg13g2_decap_8
XFILLER_15_56 VPWR VGND sg13g2_decap_8
XFILLER_40_147 VPWR VGND sg13g2_decap_8
X_09317_ _03469_ VPWR _03470_ VGND _03394_ _03392_ sg13g2_o21ai_1
XFILLER_15_67 VPWR VGND sg13g2_fill_2
XFILLER_22_862 VPWR VGND sg13g2_decap_4
XFILLER_22_884 VPWR VGND sg13g2_decap_8
X_09248_ _03399_ _03401_ _03402_ VPWR VGND sg13g2_nor2_1
Xclkbuf_4_10_0_clk clknet_0_clk clknet_4_10_0_clk VPWR VGND sg13g2_buf_8
XFILLER_108_923 VPWR VGND sg13g2_decap_8
X_09179_ _03342_ VPWR _01287_ VGND net1899 _03341_ sg13g2_o21ai_1
XFILLER_5_527 VPWR VGND sg13g2_decap_8
XFILLER_31_77 VPWR VGND sg13g2_decap_4
XFILLER_123_904 VPWR VGND sg13g2_decap_8
X_11210_ _05121_ _05111_ _05130_ _05176_ VPWR VGND sg13g2_nand3_1
X_12190_ _06036_ _06030_ _06035_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_88 VPWR VGND sg13g2_decap_8
XFILLER_31_99 VPWR VGND sg13g2_fill_2
X_11141_ _05023_ _05110_ _05111_ VPWR VGND sg13g2_nor2_1
Xplace1790 net1788 net1790 VPWR VGND sg13g2_buf_2
XFILLER_0_210 VPWR VGND sg13g2_decap_8
X_11072_ _04993_ _05048_ _05049_ VPWR VGND sg13g2_nor2_2
XFILLER_0_232 VPWR VGND sg13g2_decap_8
X_14900_ _00701_ VGND VPWR _01420_ acc_sub.op_sign_logic0.mantisa_b\[10\] clknet_leaf_62_clk
+ sg13g2_dfrbpq_1
XFILLER_48_214 VPWR VGND sg13g2_decap_8
X_10023_ VPWR _04111_ _04110_ VGND sg13g2_inv_1
X_14831_ _00632_ VGND VPWR _01355_ fpdiv.divider0.remainder_reg\[10\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_2
XFILLER_76_556 VPWR VGND sg13g2_decap_8
XFILLER_56_30 VPWR VGND sg13g2_fill_1
X_14762_ _00563_ VGND VPWR _01286_ acc_sum.exp_mant_logic0.b\[7\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_11974_ _05828_ fpmul.reg_a_out\[11\] fpmul.reg_b_out\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_16_100 VPWR VGND sg13g2_fill_2
XFILLER_16_122 VPWR VGND sg13g2_fill_1
XFILLER_72_773 VPWR VGND sg13g2_fill_1
XFILLER_60_924 VPWR VGND sg13g2_fill_2
XFILLER_60_902 VPWR VGND sg13g2_decap_8
X_13713_ VPWR _00264_ net60 VGND sg13g2_inv_1
X_14693_ _00494_ VGND VPWR _01221_ fp16_res_pipe.op_sign_logic0.add_sub clknet_leaf_130_clk
+ sg13g2_dfrbpq_2
X_10925_ _04741_ VPWR _04933_ VGND _04811_ _04932_ sg13g2_o21ai_1
XFILLER_112_91 VPWR VGND sg13g2_decap_8
XFILLER_108_1007 VPWR VGND sg13g2_decap_8
XFILLER_71_272 VPWR VGND sg13g2_decap_8
X_13644_ VPWR _00195_ net111 VGND sg13g2_inv_1
XFILLER_60_946 VPWR VGND sg13g2_decap_8
X_10856_ net1824 fp16_res_pipe.add_renorm0.exp\[2\] _04868_ VPWR VGND sg13g2_nor2_1
XFILLER_31_136 VPWR VGND sg13g2_fill_2
X_13575_ VPWR _00126_ net32 VGND sg13g2_inv_1
XFILLER_13_884 VPWR VGND sg13g2_decap_8
X_10787_ _04799_ fp16_res_pipe.add_renorm0.exp\[3\] _04777_ VPWR VGND sg13g2_xnor2_1
X_12526_ _06349_ acc_sub.x2\[4\] net1955 VPWR VGND sg13g2_nand2_1
X_12457_ VGND VPWR _06299_ net1870 _00967_ _06300_ sg13g2_a21oi_1
XFILLER_9_899 VPWR VGND sg13g2_decap_8
XFILLER_126_764 VPWR VGND sg13g2_decap_8
X_11408_ _05349_ VPWR _01065_ VGND _05348_ net1706 sg13g2_o21ai_1
XFILLER_125_252 VPWR VGND sg13g2_decap_8
XFILLER_114_937 VPWR VGND sg13g2_decap_8
XFILLER_98_103 VPWR VGND sg13g2_decap_8
X_14127_ VPWR _00678_ net129 VGND sg13g2_inv_1
X_12388_ VPWR _06234_ _06233_ VGND sg13g2_inv_1
XFILLER_28_1008 VPWR VGND sg13g2_decap_4
X_11339_ _05293_ net1811 net1653 acc_sum.exp_mant_logic0.b\[4\] net1654 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_98_169 VPWR VGND sg13g2_decap_8
XFILLER_97_92 VPWR VGND sg13g2_fill_1
X_14058_ VPWR _00609_ net80 VGND sg13g2_inv_1
XFILLER_79_361 VPWR VGND sg13g2_fill_1
XFILLER_79_350 VPWR VGND sg13g2_fill_2
XFILLER_95_821 VPWR VGND sg13g2_fill_2
X_13009_ _06777_ _06776_ VPWR VGND _06775_ sg13g2_nand2b_2
XFILLER_95_854 VPWR VGND sg13g2_decap_4
XFILLER_94_342 VPWR VGND sg13g2_decap_8
XFILLER_67_589 VPWR VGND sg13g2_fill_2
XFILLER_54_217 VPWR VGND sg13g2_decap_8
X_08550_ _02771_ _02773_ _02774_ VPWR VGND sg13g2_nor2_2
X_08481_ _02710_ _02666_ _02660_ VPWR VGND sg13g2_nand2_1
X_07501_ _01439_ _01782_ _01823_ net1782 _01778_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_976 VPWR VGND sg13g2_decap_8
XFILLER_35_453 VPWR VGND sg13g2_decap_8
X_07432_ fpdiv.divider0.divisor_reg\[9\] net1749 _01765_ VPWR VGND sg13g2_nor2_1
XFILLER_62_261 VPWR VGND sg13g2_decap_8
XFILLER_51_935 VPWR VGND sg13g2_fill_2
XFILLER_35_497 VPWR VGND sg13g2_decap_8
XFILLER_50_467 VPWR VGND sg13g2_fill_1
X_09102_ VGND VPWR _03177_ _03178_ _03284_ _03206_ sg13g2_a21oi_1
X_07363_ _01718_ net1799 acc_sub.seg_reg0.q\[25\] VPWR VGND sg13g2_nand2_1
X_07294_ _01661_ _01521_ _01660_ VPWR VGND sg13g2_xnor2_1
X_09033_ net1790 _03154_ _03218_ _03219_ VPWR VGND sg13g2_a21o_1
XFILLER_11_1001 VPWR VGND sg13g2_decap_8
XFILLER_11_1012 VPWR VGND sg13g2_fill_2
XFILLER_117_753 VPWR VGND sg13g2_decap_8
XFILLER_117_14 VPWR VGND sg13g2_decap_8
XFILLER_105_937 VPWR VGND sg13g2_decap_8
XFILLER_104_436 VPWR VGND sg13g2_decap_4
XFILLER_89_114 VPWR VGND sg13g2_fill_1
XFILLER_120_918 VPWR VGND sg13g2_decap_8
XFILLER_113_970 VPWR VGND sg13g2_decap_8
X_09935_ _01220_ _03991_ _04031_ net1765 _03987_ VPWR VGND sg13g2_a22oi_1
X_09866_ net1820 acc_sum.y\[5\] _03973_ VPWR VGND sg13g2_nor2_1
XFILLER_98_692 VPWR VGND sg13g2_fill_1
XFILLER_86_821 VPWR VGND sg13g2_fill_2
X_08817_ _03004_ _03002_ _03003_ VPWR VGND sg13g2_xnor2_1
XFILLER_100_653 VPWR VGND sg13g2_fill_1
XFILLER_86_865 VPWR VGND sg13g2_fill_1
X_09797_ _03906_ _03910_ _03911_ VPWR VGND sg13g2_nor2_1
XFILLER_73_526 VPWR VGND sg13g2_decap_8
XFILLER_46_729 VPWR VGND sg13g2_decap_8
X_08748_ VPWR _02945_ acc_sum.exp_mant_logic0.a\[9\] VGND sg13g2_inv_1
XFILLER_27_932 VPWR VGND sg13g2_decap_8
X_08679_ VPWR _02895_ _02826_ VGND sg13g2_inv_1
XFILLER_53_272 VPWR VGND sg13g2_fill_1
XFILLER_53_261 VPWR VGND sg13g2_decap_8
XFILLER_42_957 VPWR VGND sg13g2_decap_8
XFILLER_42_946 VPWR VGND sg13g2_fill_1
X_10710_ _04681_ _04675_ _04723_ VPWR VGND sg13g2_nor2_1
XFILLER_26_77 VPWR VGND sg13g2_decap_8
XFILLER_41_434 VPWR VGND sg13g2_decap_8
XFILLER_13_125 VPWR VGND sg13g2_decap_8
X_11690_ _05593_ _05576_ _05594_ VPWR VGND sg13g2_nor2b_1
XFILLER_42_21 VPWR VGND sg13g2_decap_8
X_10641_ _04654_ _04652_ _04653_ VPWR VGND sg13g2_nand2_2
XFILLER_10_821 VPWR VGND sg13g2_decap_8
XFILLER_13_169 VPWR VGND sg13g2_fill_1
XFILLER_127_506 VPWR VGND sg13g2_decap_8
X_13360_ _07054_ _07027_ fp16_res_pipe.x2\[0\] VPWR VGND sg13g2_nand2_1
X_10572_ _04599_ acc_sub.x2\[13\] net1931 VPWR VGND sg13g2_nand2_1
X_13291_ acc\[5\] _07005_ net1679 _00839_ VPWR VGND sg13g2_mux2_1
X_12311_ _06157_ _06156_ _06086_ VPWR VGND sg13g2_nand2_1
XFILLER_42_98 VPWR VGND sg13g2_decap_8
XFILLER_6_836 VPWR VGND sg13g2_decap_8
XFILLER_108_731 VPWR VGND sg13g2_decap_8
XFILLER_107_230 VPWR VGND sg13g2_decap_8
X_12242_ _06088_ _06086_ _06087_ VPWR VGND sg13g2_nand2_1
XFILLER_10_898 VPWR VGND sg13g2_decap_8
XFILLER_101_0 VPWR VGND sg13g2_decap_8
X_12173_ _06013_ _06016_ _06011_ _06019_ VPWR VGND sg13g2_nand3_1
XFILLER_123_778 VPWR VGND sg13g2_decap_8
XFILLER_122_266 VPWR VGND sg13g2_decap_8
XFILLER_111_929 VPWR VGND sg13g2_decap_8
X_11124_ _05093_ VPWR _05094_ VGND _05048_ _05088_ sg13g2_o21ai_1
XFILLER_1_541 VPWR VGND sg13g2_decap_4
XFILLER_114_1000 VPWR VGND sg13g2_decap_8
XFILLER_110_428 VPWR VGND sg13g2_fill_1
XFILLER_107_91 VPWR VGND sg13g2_decap_8
XFILLER_104_992 VPWR VGND sg13g2_decap_8
X_11055_ VPWR _05033_ _05012_ VGND sg13g2_inv_1
XFILLER_77_876 VPWR VGND sg13g2_decap_8
XFILLER_67_62 VPWR VGND sg13g2_fill_2
X_10006_ _04003_ _04087_ _04094_ VPWR VGND sg13g2_nor2_1
XFILLER_76_375 VPWR VGND sg13g2_decap_4
XFILLER_37_718 VPWR VGND sg13g2_fill_1
X_14814_ _00615_ VGND VPWR _01338_ acc_sum.add_renorm0.mantisa\[3\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_83_61 VPWR VGND sg13g2_fill_1
X_11957_ VPWR _05815_ fpmul.seg_reg0.q\[27\] VGND sg13g2_inv_1
X_14745_ _00546_ VGND VPWR _01273_ fp16_res_pipe.add_renorm0.mantisa\[8\] clknet_leaf_136_clk
+ sg13g2_dfrbpq_1
XFILLER_17_453 VPWR VGND sg13g2_decap_4
XFILLER_18_976 VPWR VGND sg13g2_decap_8
XFILLER_83_72 VPWR VGND sg13g2_decap_8
XFILLER_33_946 VPWR VGND sg13g2_decap_8
X_10908_ _04915_ _04916_ _04917_ VPWR VGND sg13g2_nor2_1
X_11888_ fpdiv.divider0.state _05768_ _02647_ _05775_ VPWR VGND sg13g2_nand3_1
X_14676_ _00477_ VGND VPWR _01204_ fp16_res_pipe.op_sign_logic0.mantisa_a\[2\] clknet_leaf_144_clk
+ sg13g2_dfrbpq_2
X_13627_ VPWR _00178_ net57 VGND sg13g2_inv_1
X_10839_ _04798_ _04850_ _04851_ VPWR VGND sg13g2_nor2_2
X_13558_ VPWR _00109_ net21 VGND sg13g2_inv_1
XFILLER_118_517 VPWR VGND sg13g2_decap_4
X_12509_ VPWR _06339_ acc_sub.x2\[11\] VGND sg13g2_inv_1
XFILLER_8_140 VPWR VGND sg13g2_decap_8
X_13489_ VPWR _00040_ net87 VGND sg13g2_inv_1
XFILLER_114_734 VPWR VGND sg13g2_decap_8
XFILLER_114_723 VPWR VGND sg13g2_fill_2
XFILLER_87_607 VPWR VGND sg13g2_decap_8
Xfanout119 net128 net119 VPWR VGND sg13g2_buf_2
Xfanout108 net113 net108 VPWR VGND sg13g2_buf_2
X_07981_ _02253_ VPWR _01389_ VGND _02199_ _02248_ sg13g2_o21ai_1
X_09720_ VGND VPWR _03835_ _03836_ _03815_ net1690 sg13g2_a21oi_2
XFILLER_110_962 VPWR VGND sg13g2_decap_8
XFILLER_95_651 VPWR VGND sg13g2_decap_4
XFILLER_86_139 VPWR VGND sg13g2_decap_8
XFILLER_68_876 VPWR VGND sg13g2_decap_8
XFILLER_68_854 VPWR VGND sg13g2_decap_4
XFILLER_68_843 VPWR VGND sg13g2_decap_8
XFILLER_67_342 VPWR VGND sg13g2_fill_1
X_09651_ _03768_ _03631_ _03687_ _03767_ _03645_ VPWR VGND sg13g2_a22oi_1
XFILLER_94_150 VPWR VGND sg13g2_decap_8
XFILLER_27_217 VPWR VGND sg13g2_decap_4
X_09582_ VPWR _03699_ _03698_ VGND sg13g2_inv_1
XFILLER_83_868 VPWR VGND sg13g2_fill_1
XFILLER_82_334 VPWR VGND sg13g2_decap_8
X_08602_ VPWR _02825_ _02824_ VGND sg13g2_inv_1
XFILLER_27_239 VPWR VGND sg13g2_decap_8
X_08533_ VPWR _02757_ _02756_ VGND sg13g2_inv_1
XFILLER_82_367 VPWR VGND sg13g2_decap_4
XFILLER_36_762 VPWR VGND sg13g2_fill_2
XFILLER_35_250 VPWR VGND sg13g2_decap_8
XFILLER_23_423 VPWR VGND sg13g2_fill_1
XFILLER_24_946 VPWR VGND sg13g2_decap_8
X_08464_ VGND VPWR net1647 _02695_ _02697_ _02696_ sg13g2_a21oi_1
XFILLER_50_242 VPWR VGND sg13g2_decap_8
X_07415_ _01752_ net1894 acc\[1\] VPWR VGND sg13g2_nand2_1
X_07346_ _01706_ VPWR _01477_ VGND acc_sub.reg2en.q\[0\] _01700_ sg13g2_o21ai_1
XFILLER_12_35 VPWR VGND sg13g2_decap_8
X_09016_ VPWR _03202_ _03094_ VGND sg13g2_inv_1
X_07277_ _01646_ _01645_ _01636_ VPWR VGND sg13g2_nand2_1
XFILLER_5_7 VPWR VGND sg13g2_decap_8
X_09918_ VPWR _04015_ _04014_ VGND sg13g2_inv_1
XFILLER_86_651 VPWR VGND sg13g2_fill_2
XFILLER_59_843 VPWR VGND sg13g2_fill_2
X_09849_ _03840_ _03648_ _03959_ VPWR VGND sg13g2_nor2_1
XFILLER_101_962 VPWR VGND sg13g2_decap_8
XFILLER_100_461 VPWR VGND sg13g2_decap_8
XFILLER_59_898 VPWR VGND sg13g2_decap_8
XFILLER_46_515 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_fill_1
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_74_868 VPWR VGND sg13g2_fill_1
X_12860_ VGND VPWR net1935 add_result\[9\] _06639_ net1943 sg13g2_a21oi_1
XFILLER_2_1010 VPWR VGND sg13g2_decap_4
XFILLER_37_98 VPWR VGND sg13g2_decap_8
X_11811_ _05712_ _05711_ _05604_ VPWR VGND sg13g2_nand2_1
XFILLER_33_209 VPWR VGND sg13g2_fill_2
X_14530_ _00331_ VGND VPWR _01066_ fpdiv.div_out\[5\] clknet_leaf_75_clk sg13g2_dfrbpq_1
XFILLER_57_1012 VPWR VGND sg13g2_fill_2
XFILLER_42_721 VPWR VGND sg13g2_decap_4
XFILLER_14_401 VPWR VGND sg13g2_fill_2
XFILLER_15_924 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_fill_1
XFILLER_53_42 VPWR VGND sg13g2_decap_8
X_11742_ _05645_ VPWR _05646_ VGND _05627_ _05644_ sg13g2_o21ai_1
XFILLER_14_434 VPWR VGND sg13g2_decap_4
X_14461_ _00262_ VGND VPWR _01000_ fpmul.seg_reg0.q\[46\] clknet_leaf_92_clk sg13g2_dfrbpq_1
XFILLER_41_275 VPWR VGND sg13g2_fill_2
XFILLER_30_927 VPWR VGND sg13g2_decap_8
X_11673_ _04589_ _05576_ _05577_ VPWR VGND sg13g2_nor2_1
X_14392_ _00193_ VGND VPWR _00931_ div_result\[5\] clknet_leaf_81_clk sg13g2_dfrbpq_1
X_13412_ _07085_ net1722 instr\[11\] VPWR VGND sg13g2_nand2_1
X_10624_ _04632_ _04636_ _04637_ VPWR VGND sg13g2_nor2_1
X_13343_ _07045_ net1726 fp16_res_pipe.x2\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_127_336 VPWR VGND sg13g2_decap_8
X_10555_ _04588_ VPWR _01157_ VGND net1846 _04587_ sg13g2_o21ai_1
X_13274_ _06992_ net1711 acc_sub.y\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_6_688 VPWR VGND sg13g2_fill_2
XFILLER_5_154 VPWR VGND sg13g2_decap_8
X_10486_ _04515_ net1670 net1736 _04532_ VPWR VGND sg13g2_a21o_1
X_12225_ _06070_ _06069_ _06071_ VPWR VGND sg13g2_xor2_1
XFILLER_123_553 VPWR VGND sg13g2_decap_8
XFILLER_97_905 VPWR VGND sg13g2_decap_4
X_12156_ _06002_ _05999_ _06001_ VPWR VGND sg13g2_nand2_1
XFILLER_111_715 VPWR VGND sg13g2_decap_8
XFILLER_97_949 VPWR VGND sg13g2_decap_8
X_11107_ _05077_ _02947_ acc_sum.exp_mant_logic0.b\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_38_7 VPWR VGND sg13g2_decap_8
X_12087_ _05933_ _05930_ _05932_ VPWR VGND sg13g2_nand2_1
XFILLER_76_161 VPWR VGND sg13g2_fill_1
X_11038_ _05015_ _05016_ _05017_ VPWR VGND sg13g2_nor2_1
XFILLER_37_504 VPWR VGND sg13g2_fill_1
XFILLER_77_695 VPWR VGND sg13g2_fill_1
XFILLER_64_323 VPWR VGND sg13g2_fill_2
XFILLER_37_537 VPWR VGND sg13g2_decap_4
XFILLER_37_559 VPWR VGND sg13g2_fill_2
XFILLER_73_890 VPWR VGND sg13g2_decap_8
X_12989_ VPWR _06757_ _06756_ VGND sg13g2_inv_1
X_14728_ _00529_ VGND VPWR _01256_ fp16_res_pipe.exp_mant_logic0.a\[15\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
XFILLER_71_1009 VPWR VGND sg13g2_decap_4
X_14659_ _00460_ VGND VPWR _01187_ fp16_res_pipe.exp_mant_logic0.b\[12\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_1
XFILLER_21_938 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_32_253 VPWR VGND sg13g2_decap_8
X_07200_ VPWR _01572_ _01534_ VGND sg13g2_inv_1
X_08180_ _02438_ fp16_sum_pipe.exp_mant_logic0.a\[5\] _02408_ fp16_sum_pipe.exp_mant_logic0.a\[6\]
+ _02332_ VPWR VGND sg13g2_a22oi_1
X_07131_ VPWR _01503_ acc_sub.op_sign_logic0.mantisa_a\[8\] VGND sg13g2_inv_1
XFILLER_118_336 VPWR VGND sg13g2_fill_1
XFILLER_64_0 VPWR VGND sg13g2_fill_2
XFILLER_114_564 VPWR VGND sg13g2_decap_4
XFILLER_114_586 VPWR VGND sg13g2_decap_8
XFILLER_102_715 VPWR VGND sg13g2_decap_8
XFILLER_87_437 VPWR VGND sg13g2_fill_1
XFILLER_4_91 VPWR VGND sg13g2_decap_8
X_07964_ _02238_ fp16_sum_pipe.exp_mant_logic0.a\[14\] VPWR VGND sg13g2_inv_2
X_09703_ _03799_ _03818_ _03819_ VPWR VGND sg13g2_nor2_1
X_07895_ _02174_ VPWR _01396_ VGND net1891 _02087_ sg13g2_o21ai_1
X_09634_ _03675_ _03680_ _03751_ VPWR VGND sg13g2_nor2_1
XFILLER_67_161 VPWR VGND sg13g2_decap_8
XFILLER_83_654 VPWR VGND sg13g2_decap_8
XFILLER_71_849 VPWR VGND sg13g2_fill_2
XFILLER_70_304 VPWR VGND sg13g2_fill_1
X_08516_ acc_sum.op_sign_logic0.mantisa_b\[6\] _02739_ _02740_ VPWR VGND sg13g2_nor2_2
XFILLER_24_732 VPWR VGND sg13g2_fill_1
X_09496_ _03615_ fp16_res_pipe.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_inv_2
X_08447_ VGND VPWR _02679_ _02680_ _02681_ fpdiv.divider0.divisor_reg\[11\] sg13g2_a21oi_1
XFILLER_24_787 VPWR VGND sg13g2_decap_4
XFILLER_8_909 VPWR VGND sg13g2_decap_8
XFILLER_11_426 VPWR VGND sg13g2_decap_8
X_08378_ _02619_ _02572_ _07115_ VPWR VGND sg13g2_nor2b_1
XFILLER_23_56 VPWR VGND sg13g2_decap_8
X_07329_ net1744 _01602_ _01691_ _01692_ VPWR VGND sg13g2_nand3_1
XFILLER_109_336 VPWR VGND sg13g2_fill_1
XFILLER_109_325 VPWR VGND sg13g2_decap_8
X_10340_ VPWR _04390_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[8\] VGND sg13g2_inv_1
XFILLER_105_520 VPWR VGND sg13g2_decap_8
X_10271_ _04341_ _04177_ fp16_res_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
X_12010_ VGND VPWR _05861_ net1875 _00976_ _05862_ sg13g2_a21oi_1
XFILLER_105_597 VPWR VGND sg13g2_decap_4
XFILLER_105_586 VPWR VGND sg13g2_fill_1
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_94_919 VPWR VGND sg13g2_decap_8
XFILLER_78_437 VPWR VGND sg13g2_decap_4
XFILLER_59_640 VPWR VGND sg13g2_decap_4
XFILLER_48_42 VPWR VGND sg13g2_decap_8
X_13961_ VPWR _00512_ net97 VGND sg13g2_inv_1
XFILLER_19_504 VPWR VGND sg13g2_decap_8
XFILLER_100_280 VPWR VGND sg13g2_decap_8
XFILLER_87_993 VPWR VGND sg13g2_decap_8
XFILLER_86_470 VPWR VGND sg13g2_fill_2
X_12912_ _06687_ _06683_ _06686_ _06516_ net1949 VPWR VGND sg13g2_a22oi_1
XFILLER_0_49 VPWR VGND sg13g2_decap_8
X_13892_ VPWR _00443_ net43 VGND sg13g2_inv_1
X_12843_ _06624_ _06623_ net1732 VPWR VGND sg13g2_nand2_1
XFILLER_62_827 VPWR VGND sg13g2_decap_8
XFILLER_61_315 VPWR VGND sg13g2_decap_8
XFILLER_15_721 VPWR VGND sg13g2_fill_1
XFILLER_27_570 VPWR VGND sg13g2_decap_4
X_12774_ _06556_ _06558_ _06559_ VPWR VGND sg13g2_nor2b_2
XFILLER_61_348 VPWR VGND sg13g2_decap_8
XFILLER_14_231 VPWR VGND sg13g2_decap_8
X_14513_ _00314_ VGND VPWR _01049_ fpdiv.divider0.dividend\[8\] clknet_leaf_85_clk
+ sg13g2_dfrbpq_1
X_11725_ _05629_ _05624_ _05628_ VPWR VGND sg13g2_nand2_1
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_14_242 VPWR VGND sg13g2_fill_1
XFILLER_14_264 VPWR VGND sg13g2_fill_1
XFILLER_15_787 VPWR VGND sg13g2_decap_4
XFILLER_30_713 VPWR VGND sg13g2_fill_2
XFILLER_120_91 VPWR VGND sg13g2_decap_8
X_14444_ _00245_ VGND VPWR _00983_ fpmul.seg_reg0.q\[29\] clknet_leaf_105_clk sg13g2_dfrbpq_1
Xfanout90 net91 net90 VPWR VGND sg13g2_buf_2
XFILLER_80_84 VPWR VGND sg13g2_fill_1
X_11656_ net1836 _05560_ _05561_ VPWR VGND sg13g2_nor2_1
XFILLER_30_779 VPWR VGND sg13g2_fill_2
XFILLER_127_133 VPWR VGND sg13g2_decap_8
X_14375_ _00176_ VGND VPWR _00916_ fpmul.reg_b_out\[6\] clknet_leaf_101_clk sg13g2_dfrbpq_2
X_10607_ VPWR _04620_ _04619_ VGND sg13g2_inv_1
X_11587_ _05492_ _05461_ _05484_ _05470_ VPWR VGND sg13g2_and3_1
XFILLER_116_807 VPWR VGND sg13g2_decap_8
XFILLER_109_870 VPWR VGND sg13g2_decap_4
X_13326_ _07033_ VPWR _00832_ VGND _07032_ net1725 sg13g2_o21ai_1
XFILLER_7_986 VPWR VGND sg13g2_decap_8
X_10538_ _04577_ _04474_ _04576_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_481 VPWR VGND sg13g2_decap_8
XFILLER_10_492 VPWR VGND sg13g2_fill_1
X_13257_ VGND VPWR net1679 _06978_ _00847_ _06979_ sg13g2_a21oi_1
XFILLER_6_474 VPWR VGND sg13g2_decap_8
XFILLER_124_851 VPWR VGND sg13g2_decap_8
XFILLER_89_82 VPWR VGND sg13g2_decap_8
X_12208_ VPWR _06054_ _06011_ VGND sg13g2_inv_1
X_10469_ _04505_ _04516_ _04517_ VPWR VGND sg13g2_nor2_1
X_13188_ _06926_ VPWR _00863_ VGND _06925_ net1712 sg13g2_o21ai_1
XFILLER_111_545 VPWR VGND sg13g2_decap_8
X_12139_ VGND VPWR _05923_ _05926_ _05985_ _05984_ sg13g2_a21oi_1
XFILLER_2_680 VPWR VGND sg13g2_fill_1
XFILLER_111_567 VPWR VGND sg13g2_decap_8
XFILLER_97_779 VPWR VGND sg13g2_fill_1
XFILLER_96_278 VPWR VGND sg13g2_decap_8
XFILLER_84_429 VPWR VGND sg13g2_decap_8
XFILLER_96_289 VPWR VGND sg13g2_fill_1
XFILLER_65_632 VPWR VGND sg13g2_fill_1
XFILLER_65_621 VPWR VGND sg13g2_decap_8
XFILLER_49_161 VPWR VGND sg13g2_decap_8
XFILLER_37_301 VPWR VGND sg13g2_decap_8
X_07680_ net1660 _01988_ _01989_ VPWR VGND sg13g2_nor2b_2
XFILLER_65_676 VPWR VGND sg13g2_decap_8
XFILLER_93_996 VPWR VGND sg13g2_decap_8
XFILLER_92_495 VPWR VGND sg13g2_fill_2
XFILLER_80_602 VPWR VGND sg13g2_decap_4
XFILLER_53_849 VPWR VGND sg13g2_decap_8
XFILLER_25_518 VPWR VGND sg13g2_fill_2
XFILLER_64_197 VPWR VGND sg13g2_decap_4
X_09350_ _03501_ _03447_ _03499_ _03502_ VPWR VGND sg13g2_nand3_1
XFILLER_80_679 VPWR VGND sg13g2_decap_4
X_09281_ fp16_res_pipe.op_sign_logic0.mantisa_a\[8\] _03434_ _03435_ VPWR VGND sg13g2_nor2_1
X_08301_ _02546_ _02547_ _02548_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_573 VPWR VGND sg13g2_fill_1
X_08232_ _02485_ fp16_sum_pipe.exp_mant_logic0.b\[6\] _02338_ _02275_ fp16_sum_pipe.exp_mant_logic0.b\[4\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_20_212 VPWR VGND sg13g2_decap_8
X_08163_ _02422_ net1658 fp16_sum_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_119_689 VPWR VGND sg13g2_decap_8
XFILLER_118_133 VPWR VGND sg13g2_decap_8
X_08094_ _02359_ net1691 fp16_sum_pipe.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_106_317 VPWR VGND sg13g2_decap_8
Xclkload71 clkload71/Y clknet_leaf_24_clk VPWR VGND sg13g2_inv_2
Xclkload60 clknet_leaf_103_clk clkload60/X VPWR VGND sg13g2_buf_8
XFILLER_115_851 VPWR VGND sg13g2_decap_8
Xclkload82 clknet_leaf_48_clk clkload82/Y VPWR VGND sg13g2_inv_4
Xclkload93 clknet_leaf_90_clk clkload93/Y VPWR VGND sg13g2_inv_4
XFILLER_47_1011 VPWR VGND sg13g2_fill_2
XFILLER_125_14 VPWR VGND sg13g2_decap_8
XFILLER_102_512 VPWR VGND sg13g2_fill_2
XFILLER_0_606 VPWR VGND sg13g2_decap_8
X_08996_ _03181_ _03145_ _03182_ VPWR VGND sg13g2_nor2_1
XFILLER_88_768 VPWR VGND sg13g2_decap_8
XFILLER_87_223 VPWR VGND sg13g2_decap_8
XFILLER_102_556 VPWR VGND sg13g2_fill_2
X_07947_ _02213_ _02221_ _02222_ VPWR VGND sg13g2_nor2_1
XFILLER_75_429 VPWR VGND sg13g2_decap_8
XFILLER_28_301 VPWR VGND sg13g2_decap_8
XFILLER_84_952 VPWR VGND sg13g2_decap_8
X_07878_ _02166_ net1886 acc_sub.x2\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_56_643 VPWR VGND sg13g2_decap_8
XFILLER_18_56 VPWR VGND sg13g2_decap_8
XFILLER_28_334 VPWR VGND sg13g2_decap_4
X_09617_ VPWR _03734_ _03733_ VGND sg13g2_inv_1
XFILLER_28_389 VPWR VGND sg13g2_fill_2
X_09548_ VPWR _03665_ _03664_ VGND sg13g2_inv_1
XFILLER_70_145 VPWR VGND sg13g2_fill_2
XFILLER_43_348 VPWR VGND sg13g2_decap_8
XFILLER_71_679 VPWR VGND sg13g2_decap_4
XFILLER_70_167 VPWR VGND sg13g2_fill_2
XFILLER_52_871 VPWR VGND sg13g2_fill_1
XFILLER_12_702 VPWR VGND sg13g2_decap_8
X_09479_ net1919 fp16_res_pipe.exp_mant_logic0.a\[7\] _03604_ VPWR VGND sg13g2_nor2_1
XFILLER_34_77 VPWR VGND sg13g2_decap_8
XFILLER_11_212 VPWR VGND sg13g2_decap_8
XFILLER_12_746 VPWR VGND sg13g2_decap_8
X_11510_ VGND VPWR _04465_ fp16_sum_pipe.add_renorm0.mantisa\[3\] _05415_ _05414_
+ sg13g2_a21oi_1
Xclkbuf_leaf_144_clk clknet_5_0__leaf_clk clknet_leaf_144_clk VPWR VGND sg13g2_buf_8
X_12490_ VGND VPWR _06325_ net1872 _00960_ _06326_ sg13g2_a21oi_1
XFILLER_11_245 VPWR VGND sg13g2_decap_8
X_11441_ VPWR _05370_ fpdiv.reg_a_out\[7\] VGND sg13g2_inv_1
XFILLER_50_21 VPWR VGND sg13g2_decap_8
X_14160_ VPWR _00711_ net132 VGND sg13g2_inv_1
XFILLER_109_155 VPWR VGND sg13g2_decap_4
XFILLER_109_144 VPWR VGND sg13g2_fill_1
X_11372_ _03353_ _05148_ _05323_ VPWR VGND sg13g2_nor2_1
XFILLER_125_648 VPWR VGND sg13g2_fill_1
XFILLER_109_199 VPWR VGND sg13g2_decap_8
X_13111_ _06868_ _06796_ VPWR VGND _06777_ sg13g2_nand2b_2
XFILLER_50_98 VPWR VGND sg13g2_decap_8
XFILLER_4_923 VPWR VGND sg13g2_decap_8
X_10323_ _04379_ net1920 fp16_res_pipe.x2\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_124_147 VPWR VGND sg13g2_decap_8
X_14091_ VPWR _00642_ net40 VGND sg13g2_inv_1
XFILLER_105_350 VPWR VGND sg13g2_fill_2
X_13042_ _06761_ _06809_ _06810_ VPWR VGND sg13g2_nor2_1
XFILLER_3_455 VPWR VGND sg13g2_decap_8
X_10254_ _04321_ _04324_ _04325_ VPWR VGND sg13g2_nor2_1
XFILLER_121_854 VPWR VGND sg13g2_decap_8
XFILLER_79_768 VPWR VGND sg13g2_decap_4
XFILLER_61_1008 VPWR VGND sg13g2_decap_4
XFILLER_59_63 VPWR VGND sg13g2_decap_4
X_10185_ _01202_ _04262_ _04263_ VPWR VGND sg13g2_nand2_1
XFILLER_115_91 VPWR VGND sg13g2_decap_8
XFILLER_93_226 VPWR VGND sg13g2_decap_4
XFILLER_75_941 VPWR VGND sg13g2_decap_8
XFILLER_59_470 VPWR VGND sg13g2_decap_8
XFILLER_47_632 VPWR VGND sg13g2_decap_8
X_13944_ VPWR _00495_ net27 VGND sg13g2_inv_1
XFILLER_35_805 VPWR VGND sg13g2_decap_8
XFILLER_19_334 VPWR VGND sg13g2_fill_2
XFILLER_46_175 VPWR VGND sg13g2_fill_2
XFILLER_46_153 VPWR VGND sg13g2_decap_8
XFILLER_35_849 VPWR VGND sg13g2_fill_2
X_13875_ VPWR _00426_ net53 VGND sg13g2_inv_1
XFILLER_34_304 VPWR VGND sg13g2_decap_8
XFILLER_19_389 VPWR VGND sg13g2_decap_8
X_12826_ _06608_ _06607_ _06606_ VPWR VGND sg13g2_nand2b_1
XFILLER_61_123 VPWR VGND sg13g2_decap_4
XFILLER_91_50 VPWR VGND sg13g2_fill_2
XFILLER_90_988 VPWR VGND sg13g2_decap_8
X_12757_ _06545_ fp16_res_pipe.x2\[2\] net1957 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_135_clk clknet_5_8__leaf_clk clknet_leaf_135_clk VPWR VGND sg13g2_buf_8
XFILLER_30_521 VPWR VGND sg13g2_decap_8
X_12688_ _06498_ VPWR _00935_ VGND _06496_ net1741 sg13g2_o21ai_1
X_11708_ VPWR _05612_ _05611_ VGND sg13g2_inv_1
X_14427_ _00228_ VGND VPWR _00966_ fpmul.seg_reg0.q\[12\] clknet_leaf_80_clk sg13g2_dfrbpq_1
X_11639_ _05544_ _05434_ _05494_ _05459_ _05475_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_587 VPWR VGND sg13g2_fill_2
X_14358_ _00159_ VGND VPWR _00900_ _00011_ clknet_leaf_87_clk sg13g2_dfrbpq_1
X_13309_ VPWR VGND acc_sub.y\[1\] _07019_ _02578_ net1728 _07020_ acc_sum.y\[1\] sg13g2_a221oi_1
XFILLER_115_147 VPWR VGND sg13g2_decap_8
X_14289_ _00090_ VGND VPWR _00000_ acc_sub.reg1en.d\[0\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_6_293 VPWR VGND sg13g2_decap_8
XFILLER_112_810 VPWR VGND sg13g2_decap_8
X_08850_ _03037_ net1789 acc_sub.add_renorm0.mantisa\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_112_887 VPWR VGND sg13g2_decap_8
XFILLER_111_353 VPWR VGND sg13g2_decap_8
X_07801_ _02100_ _02099_ _02063_ VPWR VGND sg13g2_nand2_1
XFILLER_97_587 VPWR VGND sg13g2_fill_1
XFILLER_97_576 VPWR VGND sg13g2_decap_8
XFILLER_57_418 VPWR VGND sg13g2_fill_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_84_204 VPWR VGND sg13g2_fill_2
X_07732_ _02038_ acc_sub.exp_mant_logic0.a\[0\] _01949_ acc_sub.exp_mant_logic0.a\[2\]
+ _01935_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_131 VPWR VGND sg13g2_decap_8
X_07663_ _01749_ _01821_ _01973_ VPWR VGND sg13g2_nor2_1
XFILLER_93_793 VPWR VGND sg13g2_decap_8
XFILLER_52_101 VPWR VGND sg13g2_fill_2
XFILLER_1_70 VPWR VGND sg13g2_decap_8
XFILLER_26_816 VPWR VGND sg13g2_fill_1
XFILLER_26_838 VPWR VGND sg13g2_fill_2
XFILLER_52_123 VPWR VGND sg13g2_decap_8
X_09402_ net1738 _03467_ _03547_ _03548_ VPWR VGND sg13g2_nand3_1
XFILLER_111_49 VPWR VGND sg13g2_decap_8
X_07594_ _01908_ _01812_ _01907_ VPWR VGND sg13g2_xnor2_1
XFILLER_81_999 VPWR VGND sg13g2_decap_8
X_09333_ _03485_ net1770 fp16_res_pipe.add_renorm0.mantisa\[10\] VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_126_clk clknet_5_13__leaf_clk clknet_leaf_126_clk VPWR VGND sg13g2_buf_8
XFILLER_52_178 VPWR VGND sg13g2_decap_4
XFILLER_40_318 VPWR VGND sg13g2_decap_4
XFILLER_21_521 VPWR VGND sg13g2_decap_8
X_09264_ VPWR _03418_ _03399_ VGND sg13g2_inv_1
XFILLER_21_554 VPWR VGND sg13g2_decap_8
XFILLER_33_392 VPWR VGND sg13g2_fill_2
X_09195_ _03353_ acc_sum.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_inv_2
X_08215_ _02461_ _02462_ _02465_ _02471_ VGND VPWR _02470_ sg13g2_nor4_2
XFILLER_101_1013 VPWR VGND sg13g2_fill_1
X_08146_ _02405_ VPWR _02406_ VGND _02262_ net1652 sg13g2_o21ai_1
XFILLER_119_497 VPWR VGND sg13g2_decap_8
XFILLER_107_615 VPWR VGND sg13g2_decap_4
XFILLER_105_7 VPWR VGND sg13g2_decap_4
XFILLER_84_1008 VPWR VGND sg13g2_decap_4
X_08077_ _02305_ _02342_ _02343_ VPWR VGND sg13g2_nor2b_2
XFILLER_20_35 VPWR VGND sg13g2_decap_8
XFILLER_106_158 VPWR VGND sg13g2_decap_8
Xplace1961 fpmul.reg1en.d\[0\] net1961 VPWR VGND sg13g2_buf_2
Xplace1950 net1948 net1950 VPWR VGND sg13g2_buf_2
XFILLER_0_414 VPWR VGND sg13g2_decap_8
XFILLER_1_948 VPWR VGND sg13g2_decap_8
XFILLER_88_576 VPWR VGND sg13g2_fill_1
XFILLER_88_565 VPWR VGND sg13g2_decap_8
X_08979_ _03165_ acc_sub.add_renorm0.exp\[0\] _03145_ VPWR VGND sg13g2_xnor2_1
XFILLER_88_587 VPWR VGND sg13g2_fill_1
XFILLER_75_259 VPWR VGND sg13g2_fill_2
XFILLER_57_952 VPWR VGND sg13g2_decap_8
X_11990_ _05837_ _05838_ _05844_ VPWR VGND sg13g2_nor2b_1
XFILLER_29_665 VPWR VGND sg13g2_fill_2
XFILLER_90_207 VPWR VGND sg13g2_fill_2
XFILLER_45_21 VPWR VGND sg13g2_decap_8
X_10941_ _04869_ _04867_ _04948_ VPWR VGND sg13g2_nor2_1
XFILLER_29_698 VPWR VGND sg13g2_decap_8
XFILLER_83_292 VPWR VGND sg13g2_decap_4
X_13660_ VPWR _00211_ net35 VGND sg13g2_inv_1
XFILLER_44_657 VPWR VGND sg13g2_fill_1
XFILLER_43_112 VPWR VGND sg13g2_decap_8
X_12611_ VPWR _06427_ _06425_ VGND sg13g2_inv_1
XFILLER_72_977 VPWR VGND sg13g2_decap_8
XFILLER_45_98 VPWR VGND sg13g2_decap_8
XFILLER_44_668 VPWR VGND sg13g2_decap_8
X_10872_ _01135_ _04882_ _04883_ VPWR VGND sg13g2_nand2_1
XFILLER_16_359 VPWR VGND sg13g2_decap_8
X_13591_ VPWR _00142_ net120 VGND sg13g2_inv_1
XFILLER_12_521 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_117_clk clknet_5_9__leaf_clk clknet_leaf_117_clk VPWR VGND sg13g2_buf_8
XFILLER_25_882 VPWR VGND sg13g2_decap_8
X_12542_ _06359_ _06357_ _06358_ VPWR VGND sg13g2_nand2_2
XFILLER_12_554 VPWR VGND sg13g2_fill_1
X_12473_ _06305_ _06146_ _06306_ _06314_ VPWR VGND sg13g2_nand3_1
XFILLER_61_75 VPWR VGND sg13g2_fill_1
X_14212_ VPWR _00763_ net135 VGND sg13g2_inv_1
X_11424_ _05359_ acc_sub.x2\[13\] VPWR VGND sg13g2_inv_2
XFILLER_126_946 VPWR VGND sg13g2_decap_8
XFILLER_125_401 VPWR VGND sg13g2_decap_4
X_14143_ VPWR _00694_ net129 VGND sg13g2_inv_1
X_11355_ _05308_ acc_sum.exp_mant_logic0.b\[0\] net1681 acc_sum.op_sign_logic0.mantisa_b\[3\]
+ net1762 VPWR VGND sg13g2_a22oi_1
XFILLER_113_618 VPWR VGND sg13g2_fill_1
XFILLER_113_607 VPWR VGND sg13g2_decap_8
XFILLER_98_318 VPWR VGND sg13g2_decap_8
X_14074_ VPWR _00625_ net94 VGND sg13g2_inv_1
X_11286_ _05247_ net1761 acc_sum.op_sign_logic0.mantisa_a\[0\] VPWR VGND sg13g2_nand2_1
X_10306_ _04370_ VPWR _01188_ VGND net1915 _04000_ sg13g2_o21ai_1
XFILLER_79_532 VPWR VGND sg13g2_fill_2
X_13025_ _06793_ net1853 fpmul.seg_reg0.q\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_4_797 VPWR VGND sg13g2_decap_8
X_10237_ _04302_ _04189_ _04309_ VPWR VGND sg13g2_nor2_1
XFILLER_39_407 VPWR VGND sg13g2_decap_8
XFILLER_121_695 VPWR VGND sg13g2_fill_1
XFILLER_120_161 VPWR VGND sg13g2_decap_8
XFILLER_94_513 VPWR VGND sg13g2_decap_8
XFILLER_86_83 VPWR VGND sg13g2_fill_1
XFILLER_66_226 VPWR VGND sg13g2_fill_1
XFILLER_20_7 VPWR VGND sg13g2_decap_8
X_10168_ _03613_ _04175_ _04248_ VPWR VGND sg13g2_nor2_1
XFILLER_94_557 VPWR VGND sg13g2_fill_2
XFILLER_82_719 VPWR VGND sg13g2_decap_8
XFILLER_82_708 VPWR VGND sg13g2_fill_1
XFILLER_48_941 VPWR VGND sg13g2_decap_4
XFILLER_19_120 VPWR VGND sg13g2_decap_8
X_10099_ _03609_ _04156_ _04183_ VPWR VGND sg13g2_nor2_1
XFILLER_75_771 VPWR VGND sg13g2_decap_8
XFILLER_63_922 VPWR VGND sg13g2_fill_2
XFILLER_35_613 VPWR VGND sg13g2_fill_2
X_13927_ VPWR _00478_ net8 VGND sg13g2_inv_1
XFILLER_63_955 VPWR VGND sg13g2_decap_8
XFILLER_35_646 VPWR VGND sg13g2_decap_8
XFILLER_34_112 VPWR VGND sg13g2_decap_8
XFILLER_90_763 VPWR VGND sg13g2_decap_4
XFILLER_63_988 VPWR VGND sg13g2_decap_8
X_13858_ VPWR _00409_ net43 VGND sg13g2_inv_1
XFILLER_23_819 VPWR VGND sg13g2_decap_4
X_12809_ _00019_ net1730 net1701 _06592_ VPWR VGND sg13g2_nand3_1
X_13789_ VPWR _00340_ net74 VGND sg13g2_inv_1
XFILLER_50_649 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_108_clk clknet_5_10__leaf_clk clknet_leaf_108_clk VPWR VGND sg13g2_buf_8
XFILLER_15_370 VPWR VGND sg13g2_decap_4
XFILLER_16_882 VPWR VGND sg13g2_decap_8
XFILLER_15_392 VPWR VGND sg13g2_fill_2
XFILLER_30_340 VPWR VGND sg13g2_fill_2
XFILLER_31_841 VPWR VGND sg13g2_decap_4
X_08000_ _02267_ fp16_sum_pipe.exp_mant_logic0.a\[6\] VPWR VGND sg13g2_inv_2
XFILLER_117_935 VPWR VGND sg13g2_decap_8
X_09951_ _04047_ _04040_ _04046_ VPWR VGND sg13g2_nand2_2
X_08902_ _03087_ _03088_ _03086_ _03089_ VPWR VGND sg13g2_nand3_1
XFILLER_97_340 VPWR VGND sg13g2_fill_1
X_09882_ _03983_ fp16_res_pipe.reg1en.d\[0\] VPWR VGND sg13g2_inv_2
X_08833_ _03020_ net1788 acc_sub.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_58_749 VPWR VGND sg13g2_decap_8
XFILLER_57_215 VPWR VGND sg13g2_fill_2
X_08764_ _02956_ acc\[4\] net1897 VPWR VGND sg13g2_nand2_1
X_07715_ _02022_ _01949_ acc_sub.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_73_719 VPWR VGND sg13g2_decap_8
XFILLER_54_922 VPWR VGND sg13g2_decap_4
X_08695_ VGND VPWR net1671 _02845_ _02909_ net1739 sg13g2_a21oi_1
XFILLER_81_730 VPWR VGND sg13g2_decap_8
XFILLER_65_292 VPWR VGND sg13g2_fill_2
XFILLER_54_955 VPWR VGND sg13g2_decap_4
XFILLER_25_123 VPWR VGND sg13g2_decap_4
X_07646_ _01958_ net1792 net1646 net1793 net1651 VPWR VGND sg13g2_a22oi_1
XFILLER_81_763 VPWR VGND sg13g2_decap_8
XFILLER_54_977 VPWR VGND sg13g2_fill_1
X_07577_ VGND VPWR _01890_ _01786_ _01891_ _01785_ sg13g2_a21oi_1
XFILLER_40_126 VPWR VGND sg13g2_decap_8
XFILLER_15_35 VPWR VGND sg13g2_decap_8
XFILLER_25_189 VPWR VGND sg13g2_fill_2
X_09316_ _03469_ _03468_ _03397_ VPWR VGND sg13g2_nand2_1
X_09247_ fp16_res_pipe.op_sign_logic0.mantisa_b\[3\] _03400_ _03401_ VPWR VGND sg13g2_nor2_1
XFILLER_21_362 VPWR VGND sg13g2_decap_8
XFILLER_108_902 VPWR VGND sg13g2_decap_8
XFILLER_21_384 VPWR VGND sg13g2_fill_2
X_09178_ _03342_ acc_sub.x2\[8\] net1897 VPWR VGND sg13g2_nand2_1
XFILLER_5_506 VPWR VGND sg13g2_decap_8
XFILLER_31_56 VPWR VGND sg13g2_decap_8
XFILLER_108_979 VPWR VGND sg13g2_decap_8
X_08129_ _02391_ fp16_sum_pipe.exp_mant_logic0.a\[2\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[5\]
+ net1776 VPWR VGND sg13g2_a22oi_1
X_11140_ _05110_ _05019_ _05109_ VPWR VGND sg13g2_xnor2_1
XFILLER_122_437 VPWR VGND sg13g2_fill_1
Xplace1780 net1779 net1780 VPWR VGND sg13g2_buf_2
Xplace1791 net1790 net1791 VPWR VGND sg13g2_buf_2
X_11071_ _05048_ _05046_ VPWR VGND sg13g2_inv_2
XFILLER_102_172 VPWR VGND sg13g2_decap_8
X_10022_ _04016_ _04109_ _04110_ VPWR VGND sg13g2_nor2_1
X_14830_ _00631_ VGND VPWR _01354_ fpdiv.divider0.remainder_reg\[9\] clknet_leaf_70_clk
+ sg13g2_dfrbpq_2
XFILLER_0_299 VPWR VGND sg13g2_decap_8
XFILLER_91_516 VPWR VGND sg13g2_decap_4
XFILLER_45_900 VPWR VGND sg13g2_fill_1
XFILLER_17_613 VPWR VGND sg13g2_decap_4
XFILLER_56_281 VPWR VGND sg13g2_decap_4
X_14761_ _00562_ VGND VPWR _01285_ acc_sum.exp_mant_logic0.b\[6\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
X_11973_ VPWR _05827_ _05826_ VGND sg13g2_inv_1
XFILLER_45_955 VPWR VGND sg13g2_decap_8
XFILLER_44_421 VPWR VGND sg13g2_fill_2
XFILLER_29_495 VPWR VGND sg13g2_fill_1
XFILLER_112_70 VPWR VGND sg13g2_decap_8
XFILLER_71_251 VPWR VGND sg13g2_decap_8
X_13712_ VPWR _00263_ net58 VGND sg13g2_inv_1
XFILLER_45_966 VPWR VGND sg13g2_fill_1
X_14692_ _00493_ VGND VPWR _01220_ fp16_res_pipe.seg_reg0.q\[29\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
X_10924_ VGND VPWR _04809_ _04740_ _04932_ _04849_ sg13g2_a21oi_1
XFILLER_32_605 VPWR VGND sg13g2_decap_8
X_13643_ VPWR _00194_ net123 VGND sg13g2_inv_1
XFILLER_72_41 VPWR VGND sg13g2_fill_2
XFILLER_60_936 VPWR VGND sg13g2_decap_8
XFILLER_16_167 VPWR VGND sg13g2_fill_1
X_10855_ _03586_ _04866_ _04867_ VPWR VGND sg13g2_nor2_1
XFILLER_32_616 VPWR VGND sg13g2_decap_4
XFILLER_32_638 VPWR VGND sg13g2_fill_2
X_13574_ VPWR _00125_ net32 VGND sg13g2_inv_1
XFILLER_13_863 VPWR VGND sg13g2_decap_8
XFILLER_25_690 VPWR VGND sg13g2_fill_2
X_12525_ _06348_ VPWR _00947_ VGND net1956 _05781_ sg13g2_o21ai_1
XFILLER_8_311 VPWR VGND sg13g2_fill_1
XFILLER_8_300 VPWR VGND sg13g2_fill_1
X_10786_ VPWR _04798_ _04797_ VGND sg13g2_inv_1
XFILLER_40_693 VPWR VGND sg13g2_decap_4
XFILLER_8_355 VPWR VGND sg13g2_fill_2
XFILLER_9_878 VPWR VGND sg13g2_decap_8
X_12456_ net1870 fpmul.seg_reg0.q\[13\] _06300_ VPWR VGND sg13g2_nor2_1
XFILLER_68_7 VPWR VGND sg13g2_fill_2
XFILLER_8_377 VPWR VGND sg13g2_fill_2
XFILLER_126_743 VPWR VGND sg13g2_decap_8
XFILLER_125_231 VPWR VGND sg13g2_decap_8
X_11407_ _05349_ net1707 fpdiv.div_out\[4\] VPWR VGND sg13g2_nand2_1
X_12387_ _06230_ _06232_ _06233_ VPWR VGND sg13g2_nor2_2
XFILLER_114_916 VPWR VGND sg13g2_decap_8
X_14126_ VPWR _00677_ net117 VGND sg13g2_inv_1
X_11338_ _05292_ acc_sum.exp_mant_logic0.b\[2\] _05161_ net1697 acc_sum.exp_mant_logic0.b\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_14057_ VPWR _00608_ net78 VGND sg13g2_inv_1
X_11269_ _05232_ net1761 acc_sum.op_sign_logic0.mantisa_a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_79_373 VPWR VGND sg13g2_decap_8
X_13008_ _06776_ net1853 fpmul.seg_reg0.q\[8\] VPWR VGND sg13g2_nand2b_1
XFILLER_121_481 VPWR VGND sg13g2_decap_4
XFILLER_79_395 VPWR VGND sg13g2_decap_8
XFILLER_82_505 VPWR VGND sg13g2_fill_2
X_14959_ _00760_ VGND VPWR _01479_ acc_sub.add_renorm0.mantisa\[3\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_2
X_07500_ _01823_ _01821_ acc_sub.exp_mant_logic0.a\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_82_549 VPWR VGND sg13g2_decap_8
XFILLER_75_590 VPWR VGND sg13g2_decap_8
XFILLER_63_741 VPWR VGND sg13g2_decap_4
XFILLER_48_793 VPWR VGND sg13g2_decap_4
XFILLER_36_955 VPWR VGND sg13g2_decap_8
X_08480_ _02709_ VPWR _01353_ VGND net1705 _02708_ sg13g2_o21ai_1
XFILLER_62_240 VPWR VGND sg13g2_decap_8
XFILLER_35_476 VPWR VGND sg13g2_decap_8
XFILLER_23_627 VPWR VGND sg13g2_decap_8
X_07362_ VPWR _01717_ acc_sub.add_renorm0.exp\[3\] VGND sg13g2_inv_1
XFILLER_94_0 VPWR VGND sg13g2_decap_8
X_09101_ _03283_ acc_sub.y\[10\] VPWR VGND sg13g2_inv_2
XFILLER_31_660 VPWR VGND sg13g2_fill_1
X_07293_ _01659_ VPWR _01660_ VGND net1667 _01657_ sg13g2_o21ai_1
X_09032_ net1790 _01717_ _03218_ VPWR VGND sg13g2_nor2_1
XFILLER_117_732 VPWR VGND sg13g2_decap_8
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_116_264 VPWR VGND sg13g2_decap_8
XFILLER_105_916 VPWR VGND sg13g2_decap_8
XFILLER_89_126 VPWR VGND sg13g2_decap_4
XFILLER_86_800 VPWR VGND sg13g2_decap_8
X_09934_ _04031_ net1703 fp16_res_pipe.exp_mant_logic0.a\[14\] VPWR VGND sg13g2_nand2_1
X_09865_ _03972_ VPWR _01231_ VGND net1768 _03775_ sg13g2_o21ai_1
XFILLER_98_682 VPWR VGND sg13g2_fill_2
X_08816_ _02966_ acc_sub.add_renorm0.mantisa\[4\] _03003_ VPWR VGND sg13g2_nor2b_1
XFILLER_100_643 VPWR VGND sg13g2_decap_4
X_09796_ VPWR _03910_ _03909_ VGND sg13g2_inv_1
XFILLER_100_676 VPWR VGND sg13g2_fill_2
XFILLER_58_579 VPWR VGND sg13g2_fill_2
XFILLER_45_218 VPWR VGND sg13g2_decap_4
XFILLER_27_911 VPWR VGND sg13g2_decap_8
XFILLER_100_698 VPWR VGND sg13g2_fill_2
X_08747_ _02944_ VPWR _01321_ VGND net1900 _02943_ sg13g2_o21ai_1
XFILLER_39_782 VPWR VGND sg13g2_decap_8
X_08678_ VGND VPWR _02893_ net1816 _01340_ _02894_ sg13g2_a21oi_1
XFILLER_53_240 VPWR VGND sg13g2_decap_8
XFILLER_26_56 VPWR VGND sg13g2_decap_8
XFILLER_27_988 VPWR VGND sg13g2_decap_8
X_07629_ _01935_ _01942_ _01943_ VPWR VGND sg13g2_nor2_1
XFILLER_81_560 VPWR VGND sg13g2_decap_4
XFILLER_54_796 VPWR VGND sg13g2_decap_8
XFILLER_13_104 VPWR VGND sg13g2_decap_8
X_10640_ VPWR _04653_ fp16_res_pipe.add_renorm0.mantisa\[10\] VGND sg13g2_inv_1
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_10_800 VPWR VGND sg13g2_decap_8
XFILLER_42_77 VPWR VGND sg13g2_decap_8
X_10571_ _04598_ VPWR _01151_ VGND net1925 _02238_ sg13g2_o21ai_1
XFILLER_108_710 VPWR VGND sg13g2_decap_8
X_13290_ _07004_ VPWR _07005_ VGND _07003_ _06952_ sg13g2_o21ai_1
X_12310_ _06156_ _06154_ _06155_ VPWR VGND sg13g2_nand2_1
XFILLER_10_877 VPWR VGND sg13g2_decap_8
X_12241_ _06087_ _06068_ _06076_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_336 VPWR VGND sg13g2_decap_8
XFILLER_108_798 VPWR VGND sg13g2_decap_4
X_12172_ _06018_ _06014_ _06017_ VPWR VGND sg13g2_nand2_1
XFILLER_1_520 VPWR VGND sg13g2_decap_8
XFILLER_123_757 VPWR VGND sg13g2_decap_8
XFILLER_122_245 VPWR VGND sg13g2_decap_8
XFILLER_111_908 VPWR VGND sg13g2_decap_8
X_11123_ _05093_ _05092_ _05026_ VPWR VGND sg13g2_nand2_1
XFILLER_104_971 VPWR VGND sg13g2_decap_8
XFILLER_89_671 VPWR VGND sg13g2_fill_1
X_11054_ VGND VPWR _05030_ _05031_ _05032_ _05015_ sg13g2_a21oi_1
XFILLER_67_30 VPWR VGND sg13g2_fill_1
XFILLER_3_49 VPWR VGND sg13g2_decap_8
X_10005_ _04092_ _04029_ _04093_ VPWR VGND _04091_ sg13g2_nand3b_1
X_14813_ _00614_ VGND VPWR _01337_ acc_sum.add_renorm0.mantisa\[2\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_76_398 VPWR VGND sg13g2_fill_2
XFILLER_76_387 VPWR VGND sg13g2_decap_8
XFILLER_18_955 VPWR VGND sg13g2_decap_8
XFILLER_123_91 VPWR VGND sg13g2_decap_8
XFILLER_91_379 VPWR VGND sg13g2_fill_2
XFILLER_91_368 VPWR VGND sg13g2_decap_8
X_11956_ _05814_ VPWR _00982_ VGND net1883 _05813_ sg13g2_o21ai_1
X_14744_ _00545_ VGND VPWR _01272_ fp16_res_pipe.add_renorm0.mantisa\[7\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_2
XFILLER_17_432 VPWR VGND sg13g2_decap_8
XFILLER_44_262 VPWR VGND sg13g2_fill_1
XFILLER_44_251 VPWR VGND sg13g2_fill_2
XFILLER_33_925 VPWR VGND sg13g2_decap_8
X_10907_ VPWR _04916_ _04850_ VGND sg13g2_inv_1
X_11887_ VPWR _05774_ fpdiv.divider0.counter\[1\] VGND sg13g2_inv_1
XFILLER_60_766 VPWR VGND sg13g2_decap_4
X_14675_ _00476_ VGND VPWR _01203_ fp16_res_pipe.op_sign_logic0.mantisa_a\[1\] clknet_leaf_144_clk
+ sg13g2_dfrbpq_2
X_13626_ VPWR _00177_ net61 VGND sg13g2_inv_1
XFILLER_9_620 VPWR VGND sg13g2_decap_8
XFILLER_20_608 VPWR VGND sg13g2_fill_2
X_10838_ _04850_ _04848_ _04849_ VPWR VGND sg13g2_nand2_2
X_13557_ VPWR _00108_ net21 VGND sg13g2_inv_1
X_10769_ _04781_ _04780_ fp16_res_pipe.add_renorm0.exp\[6\] VPWR VGND sg13g2_nand2_1
X_13488_ VPWR _00039_ net83 VGND sg13g2_inv_1
X_12508_ VGND VPWR _06337_ net1953 _00954_ _06338_ sg13g2_a21oi_1
X_12439_ _06272_ _06284_ _06285_ VPWR VGND sg13g2_nor2b_1
XFILLER_8_196 VPWR VGND sg13g2_decap_8
XFILLER_126_540 VPWR VGND sg13g2_decap_4
XFILLER_114_702 VPWR VGND sg13g2_fill_1
XFILLER_99_402 VPWR VGND sg13g2_fill_1
XFILLER_113_223 VPWR VGND sg13g2_decap_4
XFILLER_5_892 VPWR VGND sg13g2_decap_8
Xfanout109 net113 net109 VPWR VGND sg13g2_buf_1
X_07980_ _02253_ fp16_sum_pipe.exp_mant_logic0.a\[12\] _02250_ fp16_sum_pipe.seg_reg0.q\[27\]
+ net1775 VPWR VGND sg13g2_a22oi_1
X_14109_ VPWR _00660_ net46 VGND sg13g2_inv_1
XFILLER_80_1011 VPWR VGND sg13g2_fill_2
X_09650_ _03767_ _03628_ _03640_ VPWR VGND sg13g2_nand2_1
XFILLER_110_941 VPWR VGND sg13g2_decap_8
XFILLER_95_630 VPWR VGND sg13g2_decap_8
XFILLER_95_685 VPWR VGND sg13g2_decap_8
XFILLER_83_825 VPWR VGND sg13g2_decap_8
X_08601_ _02824_ acc_sum.op_sign_logic0.mantisa_a\[3\] acc_sum.op_sign_logic0.mantisa_b\[3\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_28_719 VPWR VGND sg13g2_decap_8
XFILLER_103_39 VPWR VGND sg13g2_decap_8
X_09581_ _03698_ net1805 acc_sum.add_renorm0.mantisa\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_82_324 VPWR VGND sg13g2_decap_4
X_08532_ _02748_ _02755_ _02756_ VPWR VGND sg13g2_nor2_2
X_08463_ net1647 fpdiv.divider0.remainder_reg\[10\] _02696_ VPWR VGND sg13g2_nor2b_1
XFILLER_91_880 VPWR VGND sg13g2_fill_1
XFILLER_36_785 VPWR VGND sg13g2_decap_8
XFILLER_24_925 VPWR VGND sg13g2_decap_8
X_07414_ _01751_ acc_sub.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_inv_2
XFILLER_23_457 VPWR VGND sg13g2_decap_8
X_08394_ _02631_ _02630_ _02563_ VPWR VGND sg13g2_nand2_1
XFILLER_51_777 VPWR VGND sg13g2_decap_8
X_07345_ _01705_ VPWR _01706_ VGND _01495_ _01701_ sg13g2_o21ai_1
XFILLER_50_298 VPWR VGND sg13g2_fill_2
X_07276_ _01645_ _01513_ _01644_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_30_clk clknet_5_16__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
XFILLER_12_14 VPWR VGND sg13g2_decap_8
XFILLER_31_490 VPWR VGND sg13g2_fill_2
X_09015_ _03099_ _03200_ _03201_ VPWR VGND sg13g2_nor2_1
XFILLER_88_18 VPWR VGND sg13g2_decap_8
XFILLER_117_595 VPWR VGND sg13g2_fill_1
XFILLER_2_339 VPWR VGND sg13g2_decap_8
XFILLER_104_256 VPWR VGND sg13g2_decap_8
X_09917_ _04014_ _04012_ fp16_res_pipe.exp_mant_logic0.a\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_101_941 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_97_clk clknet_5_11__leaf_clk clknet_leaf_97_clk VPWR VGND sg13g2_buf_8
X_09848_ _03958_ acc_sum.add_renorm0.exp\[1\] _03957_ VPWR VGND sg13g2_xnor2_1
XFILLER_59_877 VPWR VGND sg13g2_decap_8
XFILLER_58_376 VPWR VGND sg13g2_decap_4
X_09779_ _03894_ _03867_ _03882_ VPWR VGND sg13g2_xnor2_1
XFILLER_100_473 VPWR VGND sg13g2_decap_8
XFILLER_85_184 VPWR VGND sg13g2_decap_8
XFILLER_73_335 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
X_11810_ _05711_ _05620_ _05592_ VPWR VGND sg13g2_nand2_1
XFILLER_15_903 VPWR VGND sg13g2_decap_8
X_11741_ VPWR _05645_ _05587_ VGND sg13g2_inv_1
XFILLER_27_796 VPWR VGND sg13g2_decap_8
XFILLER_53_21 VPWR VGND sg13g2_decap_8
XFILLER_30_906 VPWR VGND sg13g2_decap_8
X_14460_ _00261_ VGND VPWR _00999_ fpmul.seg_reg0.q\[45\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_41_265 VPWR VGND sg13g2_decap_8
XFILLER_14_479 VPWR VGND sg13g2_fill_2
X_11672_ fp16_sum_pipe.add_renorm0.exp\[1\] fp16_sum_pipe.add_renorm0.exp\[0\] fp16_sum_pipe.add_renorm0.exp\[2\]
+ _05576_ VPWR VGND sg13g2_nand3_1
X_14391_ _00192_ VGND VPWR _00930_ div_result\[4\] clknet_leaf_81_clk sg13g2_dfrbpq_1
X_10623_ _04631_ _04635_ _04636_ VPWR VGND sg13g2_nor2_1
XFILLER_127_315 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_21_clk clknet_5_18__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
X_13342_ VPWR _07044_ sipo.word\[8\] VGND sg13g2_inv_1
X_10554_ _04588_ fp16_sum_pipe.seg_reg0.q\[26\] net1846 VPWR VGND sg13g2_nand2_1
XFILLER_22_490 VPWR VGND sg13g2_fill_1
XFILLER_108_562 VPWR VGND sg13g2_decap_8
X_13273_ VGND VPWR net1676 _06990_ _00843_ _06991_ sg13g2_a21oi_1
XFILLER_5_133 VPWR VGND sg13g2_decap_8
X_10485_ _04522_ _04530_ _04531_ VPWR VGND sg13g2_nor2_1
XFILLER_123_521 VPWR VGND sg13g2_decap_4
XFILLER_123_510 VPWR VGND sg13g2_fill_1
X_12224_ _06070_ net1859 fpmul.reg_b_out\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_123_532 VPWR VGND sg13g2_decap_8
XFILLER_118_91 VPWR VGND sg13g2_decap_8
XFILLER_78_51 VPWR VGND sg13g2_decap_8
X_12155_ _06001_ _06000_ _05989_ VPWR VGND sg13g2_nand2_1
XFILLER_97_928 VPWR VGND sg13g2_decap_8
XFILLER_68_118 VPWR VGND sg13g2_fill_1
XFILLER_2_884 VPWR VGND sg13g2_decap_8
XFILLER_110_226 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_88_clk clknet_5_24__leaf_clk clknet_leaf_88_clk VPWR VGND sg13g2_buf_8
X_12086_ _05932_ _05931_ _05907_ VPWR VGND sg13g2_nand2_1
XFILLER_1_394 VPWR VGND sg13g2_decap_8
X_11037_ acc_sum.exp_mant_logic0.a\[9\] _03339_ _05016_ VPWR VGND sg13g2_nor2_1
XFILLER_65_814 VPWR VGND sg13g2_fill_1
XFILLER_65_803 VPWR VGND sg13g2_decap_8
XFILLER_65_836 VPWR VGND sg13g2_decap_8
XFILLER_91_143 VPWR VGND sg13g2_decap_8
XFILLER_18_763 VPWR VGND sg13g2_decap_4
X_12988_ _06756_ _05863_ _06755_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_785 VPWR VGND sg13g2_fill_2
X_11939_ VPWR _05803_ fpmul.seg_reg0.q\[33\] VGND sg13g2_inv_1
X_14727_ _00528_ VGND VPWR _01255_ fp16_res_pipe.exp_mant_logic0.a\[14\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
XFILLER_33_755 VPWR VGND sg13g2_fill_2
XFILLER_33_733 VPWR VGND sg13g2_fill_1
X_14658_ _00459_ VGND VPWR _01186_ fp16_res_pipe.exp_mant_logic0.b\[11\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
XFILLER_21_917 VPWR VGND sg13g2_decap_8
X_13609_ VPWR _00160_ net111 VGND sg13g2_inv_1
XFILLER_118_304 VPWR VGND sg13g2_fill_2
X_07130_ acc_sub.op_sign_logic0.mantisa_a\[10\] _01501_ _01502_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_12_clk clknet_5_6__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_14589_ _00390_ VGND VPWR _01121_ fp16_res_pipe.y\[0\] clknet_leaf_128_clk sg13g2_dfrbpq_1
XFILLER_119_849 VPWR VGND sg13g2_decap_8
XFILLER_9_472 VPWR VGND sg13g2_decap_8
XFILLER_118_359 VPWR VGND sg13g2_decap_8
XFILLER_57_0 VPWR VGND sg13g2_decap_8
XFILLER_114_543 VPWR VGND sg13g2_decap_8
XFILLER_88_939 VPWR VGND sg13g2_decap_8
XFILLER_88_928 VPWR VGND sg13g2_decap_8
XFILLER_87_416 VPWR VGND sg13g2_decap_8
XFILLER_4_70 VPWR VGND sg13g2_decap_8
XFILLER_102_749 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_79_clk clknet_5_26__leaf_clk clknet_leaf_79_clk VPWR VGND sg13g2_buf_8
X_07963_ _02236_ VPWR _02237_ VGND _02200_ _02235_ sg13g2_o21ai_1
XFILLER_114_49 VPWR VGND sg13g2_decap_8
X_09702_ _03818_ _03813_ _03817_ VPWR VGND sg13g2_nand2_1
XFILLER_96_983 VPWR VGND sg13g2_decap_8
X_07894_ _02174_ net1891 acc_sub.x2\[2\] VPWR VGND sg13g2_nand2_1
X_09633_ _03750_ _03691_ _03716_ VPWR VGND sg13g2_xnor2_1
XFILLER_67_173 VPWR VGND sg13g2_fill_1
XFILLER_56_825 VPWR VGND sg13g2_fill_2
XFILLER_55_313 VPWR VGND sg13g2_decap_8
XFILLER_28_538 VPWR VGND sg13g2_fill_1
X_09564_ _03678_ _03680_ _03681_ VPWR VGND _03666_ sg13g2_nand3b_1
X_08515_ VPWR _02739_ acc_sum.op_sign_logic0.mantisa_a\[6\] VGND sg13g2_inv_1
XFILLER_83_688 VPWR VGND sg13g2_decap_8
XFILLER_82_176 VPWR VGND sg13g2_fill_1
XFILLER_64_880 VPWR VGND sg13g2_decap_8
XFILLER_82_198 VPWR VGND sg13g2_decap_4
XFILLER_70_349 VPWR VGND sg13g2_fill_1
XFILLER_64_891 VPWR VGND sg13g2_fill_2
XFILLER_23_221 VPWR VGND sg13g2_decap_4
X_09495_ _03614_ VPWR _01243_ VGND net1917 _03613_ sg13g2_o21ai_1
X_08446_ _02680_ _01760_ fpdiv.divider0.remainder_reg\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_24_766 VPWR VGND sg13g2_fill_1
X_08377_ _02619_ _02559_ state\[2\] VPWR VGND sg13g2_nand2_2
XFILLER_12_939 VPWR VGND sg13g2_decap_8
XFILLER_23_35 VPWR VGND sg13g2_decap_8
XFILLER_23_276 VPWR VGND sg13g2_fill_1
XFILLER_23_287 VPWR VGND sg13g2_decap_8
XFILLER_24_799 VPWR VGND sg13g2_decap_8
X_07328_ _01691_ _01558_ _01601_ VPWR VGND sg13g2_nand2b_1
XFILLER_11_449 VPWR VGND sg13g2_fill_1
XFILLER_99_28 VPWR VGND sg13g2_decap_8
XFILLER_20_983 VPWR VGND sg13g2_decap_8
X_07259_ VGND VPWR _01628_ _01572_ _01629_ _01532_ sg13g2_a21oi_1
XFILLER_124_329 VPWR VGND sg13g2_decap_8
XFILLER_117_370 VPWR VGND sg13g2_fill_1
XFILLER_3_615 VPWR VGND sg13g2_decap_8
X_10270_ _04337_ _04339_ _04340_ VPWR VGND sg13g2_nor2_1
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
X_13960_ VPWR _00511_ net96 VGND sg13g2_inv_1
XFILLER_87_972 VPWR VGND sg13g2_decap_8
X_12911_ _06685_ _06684_ net1922 _06686_ VPWR VGND sg13g2_a21o_2
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_19_538 VPWR VGND sg13g2_fill_1
XFILLER_62_806 VPWR VGND sg13g2_fill_1
XFILLER_46_357 VPWR VGND sg13g2_decap_8
X_13891_ VPWR _00442_ net53 VGND sg13g2_inv_1
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_73_176 VPWR VGND sg13g2_decap_8
X_12842_ _06622_ VPWR _06623_ VGND net1960 _06620_ sg13g2_o21ai_1
XFILLER_55_880 VPWR VGND sg13g2_decap_8
XFILLER_15_711 VPWR VGND sg13g2_fill_1
X_12773_ _06558_ _06557_ _02623_ VPWR VGND sg13g2_nand2_2
X_14512_ _00313_ VGND VPWR _01048_ fpdiv.divider0.dividend\[7\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_1
X_11724_ VPWR _05628_ _05627_ VGND sg13g2_inv_1
XFILLER_15_766 VPWR VGND sg13g2_decap_8
XFILLER_120_70 VPWR VGND sg13g2_decap_8
XFILLER_70_1010 VPWR VGND sg13g2_decap_4
X_14443_ _00244_ VGND VPWR _00982_ fpmul.seg_reg0.q\[28\] clknet_leaf_104_clk sg13g2_dfrbpq_1
XFILLER_42_585 VPWR VGND sg13g2_decap_8
XFILLER_15_799 VPWR VGND sg13g2_fill_1
X_11655_ _05560_ _05421_ _05418_ VPWR VGND sg13g2_xnor2_1
Xfanout91 net92 net91 VPWR VGND sg13g2_buf_1
Xfanout80 net81 net80 VPWR VGND sg13g2_buf_2
XFILLER_30_769 VPWR VGND sg13g2_fill_2
XFILLER_31_1005 VPWR VGND sg13g2_decap_8
XFILLER_127_112 VPWR VGND sg13g2_decap_8
X_14374_ _00175_ VGND VPWR _00915_ fpmul.reg_b_out\[5\] clknet_leaf_106_clk sg13g2_dfrbpq_2
XFILLER_11_994 VPWR VGND sg13g2_decap_8
X_10606_ VGND VPWR _04616_ fp16_res_pipe.add_renorm0.mantisa\[3\] _04619_ _04618_
+ sg13g2_a21oi_1
X_11586_ _05491_ _05490_ _05444_ VPWR VGND sg13g2_nand2_2
X_13325_ _07033_ net1725 fp16_res_pipe.x2\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_7_965 VPWR VGND sg13g2_decap_8
XFILLER_6_453 VPWR VGND sg13g2_decap_8
X_10537_ _04576_ _04574_ _04575_ _04473_ net1737 VPWR VGND sg13g2_a22oi_1
XFILLER_127_189 VPWR VGND sg13g2_decap_8
XFILLER_109_893 VPWR VGND sg13g2_decap_8
XFILLER_108_370 VPWR VGND sg13g2_decap_8
X_13256_ acc\[13\] net1679 _06979_ VPWR VGND sg13g2_nor2_1
XFILLER_50_7 VPWR VGND sg13g2_decap_8
X_10468_ VPWR VGND _04455_ _04394_ _04515_ _04452_ _04516_ _04397_ sg13g2_a221oi_1
XFILLER_124_830 VPWR VGND sg13g2_decap_8
X_12207_ _06053_ _06024_ _06052_ VPWR VGND sg13g2_xnor2_1
XFILLER_97_736 VPWR VGND sg13g2_decap_8
X_13187_ _06926_ net1712 sipo.word\[8\] VPWR VGND sg13g2_nand2_1
X_10399_ VGND VPWR _04402_ _04407_ _04449_ _04401_ sg13g2_a21oi_1
XFILLER_96_235 VPWR VGND sg13g2_decap_8
X_12138_ _05910_ _05922_ _05984_ VPWR VGND sg13g2_nor2_1
XFILLER_84_408 VPWR VGND sg13g2_decap_8
X_12069_ fpmul.reg_a_out\[2\] net1863 net1857 _05915_ VPWR VGND sg13g2_nand3_1
XFILLER_49_140 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_1_clk clknet_5_1__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
XFILLER_49_151 VPWR VGND sg13g2_fill_1
XFILLER_93_975 VPWR VGND sg13g2_decap_8
XFILLER_64_132 VPWR VGND sg13g2_decap_4
XFILLER_38_869 VPWR VGND sg13g2_decap_8
XFILLER_92_463 VPWR VGND sg13g2_fill_2
XFILLER_80_625 VPWR VGND sg13g2_fill_2
XFILLER_64_176 VPWR VGND sg13g2_fill_2
XFILLER_64_165 VPWR VGND sg13g2_fill_2
XFILLER_52_316 VPWR VGND sg13g2_decap_4
XFILLER_52_327 VPWR VGND sg13g2_decap_8
XFILLER_61_850 VPWR VGND sg13g2_decap_8
X_08300_ _02547_ net1657 fp16_sum_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
X_09280_ VPWR _03434_ fp16_res_pipe.op_sign_logic0.mantisa_b\[8\] VGND sg13g2_inv_1
X_08231_ _01370_ _02483_ _02484_ VPWR VGND sg13g2_nand2_1
XFILLER_21_725 VPWR VGND sg13g2_decap_8
XFILLER_119_602 VPWR VGND sg13g2_fill_2
XFILLER_20_246 VPWR VGND sg13g2_decap_8
XFILLER_118_112 VPWR VGND sg13g2_decap_8
X_08162_ _02420_ VPWR _02421_ VGND _02270_ net1652 sg13g2_o21ai_1
XFILLER_119_668 VPWR VGND sg13g2_fill_1
XFILLER_119_657 VPWR VGND sg13g2_decap_8
X_08093_ _02358_ net1659 _02273_ VPWR VGND sg13g2_nand2_1
XFILLER_118_189 VPWR VGND sg13g2_decap_8
XFILLER_109_49 VPWR VGND sg13g2_decap_8
Xclkload61 clknet_leaf_105_clk clkload61/X VPWR VGND sg13g2_buf_1
Xclkload50 clknet_leaf_111_clk clkload50/X VPWR VGND sg13g2_buf_8
XFILLER_115_830 VPWR VGND sg13g2_decap_8
Xclkload83 clknet_leaf_36_clk clkload83/Y VPWR VGND sg13g2_inv_4
Xclkload72 clknet_leaf_31_clk clkload72/Y VPWR VGND sg13g2_inv_4
Xclkload94 clknet_leaf_57_clk clkload94/Y VPWR VGND sg13g2_inv_4
XFILLER_88_703 VPWR VGND sg13g2_fill_1
XFILLER_87_202 VPWR VGND sg13g2_decap_8
XFILLER_114_395 VPWR VGND sg13g2_decap_8
X_08995_ _03181_ acc_sub.add_renorm0.exp\[5\] _03141_ VPWR VGND sg13g2_xnor2_1
XFILLER_102_535 VPWR VGND sg13g2_fill_1
XFILLER_87_246 VPWR VGND sg13g2_fill_1
XFILLER_75_408 VPWR VGND sg13g2_decap_8
X_07946_ _02221_ _02215_ _02220_ VPWR VGND sg13g2_nand2_2
XFILLER_84_931 VPWR VGND sg13g2_decap_8
XFILLER_18_35 VPWR VGND sg13g2_decap_8
XFILLER_95_290 VPWR VGND sg13g2_fill_1
X_07877_ _02165_ VPWR _01405_ VGND net1888 _01799_ sg13g2_o21ai_1
XFILLER_68_493 VPWR VGND sg13g2_decap_8
X_09616_ _03733_ _03731_ _03732_ VPWR VGND sg13g2_nand2_1
XFILLER_83_485 VPWR VGND sg13g2_decap_4
XFILLER_71_625 VPWR VGND sg13g2_fill_1
XFILLER_71_614 VPWR VGND sg13g2_fill_1
XFILLER_71_603 VPWR VGND sg13g2_fill_1
XFILLER_56_699 VPWR VGND sg13g2_decap_8
XFILLER_44_828 VPWR VGND sg13g2_fill_2
XFILLER_44_817 VPWR VGND sg13g2_fill_1
X_09547_ _03648_ _03663_ _03664_ VPWR VGND sg13g2_nor2_1
XFILLER_93_1010 VPWR VGND sg13g2_decap_4
XFILLER_71_658 VPWR VGND sg13g2_decap_8
XFILLER_55_198 VPWR VGND sg13g2_decap_8
XFILLER_55_187 VPWR VGND sg13g2_decap_4
XFILLER_51_382 VPWR VGND sg13g2_fill_2
X_09478_ acc_sub.x2\[7\] _03603_ VPWR VGND sg13g2_inv_4
XFILLER_34_56 VPWR VGND sg13g2_decap_8
XFILLER_24_585 VPWR VGND sg13g2_fill_2
X_08429_ VPWR _02663_ _02662_ VGND sg13g2_inv_1
X_11440_ VGND VPWR _03601_ net1940 _01053_ _05369_ sg13g2_a21oi_1
XFILLER_7_217 VPWR VGND sg13g2_decap_4
Xclkload0 clkload0/Y clknet_5_0__leaf_clk VPWR VGND sg13g2_inv_2
X_11371_ _03357_ _05173_ _05322_ VPWR VGND sg13g2_nor2_1
XFILLER_4_902 VPWR VGND sg13g2_decap_8
XFILLER_20_791 VPWR VGND sg13g2_decap_8
XFILLER_109_178 VPWR VGND sg13g2_fill_1
XFILLER_109_167 VPWR VGND sg13g2_decap_8
X_13110_ _06867_ VPWR _00882_ VGND net1862 _06699_ sg13g2_o21ai_1
XFILLER_50_77 VPWR VGND sg13g2_decap_8
X_14090_ VPWR _00641_ net40 VGND sg13g2_inv_1
X_10322_ _04378_ VPWR _01180_ VGND net1921 _04288_ sg13g2_o21ai_1
XFILLER_124_126 VPWR VGND sg13g2_decap_8
X_13041_ VPWR _06809_ _06808_ VGND sg13g2_inv_1
XFILLER_3_434 VPWR VGND sg13g2_decap_8
Xclkbuf_5_29__f_clk clknet_4_14_0_clk clknet_5_29__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_106_885 VPWR VGND sg13g2_fill_1
XFILLER_59_42 VPWR VGND sg13g2_decap_8
XFILLER_4_979 VPWR VGND sg13g2_decap_8
X_10253_ _04323_ VPWR _04324_ VGND _04322_ net1703 sg13g2_o21ai_1
XFILLER_121_833 VPWR VGND sg13g2_decap_8
X_10184_ _04263_ net1764 fp16_res_pipe.op_sign_logic0.mantisa_a\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_120_354 VPWR VGND sg13g2_fill_2
XFILLER_120_332 VPWR VGND sg13g2_decap_4
XFILLER_94_717 VPWR VGND sg13g2_decap_4
XFILLER_78_268 VPWR VGND sg13g2_decap_8
XFILLER_115_70 VPWR VGND sg13g2_decap_8
XFILLER_75_920 VPWR VGND sg13g2_decap_8
XFILLER_19_313 VPWR VGND sg13g2_decap_8
XFILLER_47_655 VPWR VGND sg13g2_fill_2
X_13943_ VPWR _00494_ net27 VGND sg13g2_inv_1
XFILLER_75_85 VPWR VGND sg13g2_decap_4
XFILLER_74_463 VPWR VGND sg13g2_decap_8
XFILLER_62_625 VPWR VGND sg13g2_fill_2
XFILLER_35_839 VPWR VGND sg13g2_fill_1
X_13874_ VPWR _00425_ net45 VGND sg13g2_inv_1
XFILLER_90_967 VPWR VGND sg13g2_decap_8
XFILLER_74_496 VPWR VGND sg13g2_fill_2
XFILLER_62_647 VPWR VGND sg13g2_fill_2
X_12825_ VGND VPWR _04902_ net1911 _06607_ net1924 sg13g2_a21oi_1
XFILLER_61_168 VPWR VGND sg13g2_fill_2
XFILLER_43_850 VPWR VGND sg13g2_fill_1
XFILLER_70_691 VPWR VGND sg13g2_decap_8
X_12756_ fpmul.reg_b_out\[3\] fp16_res_pipe.x2\[3\] net1957 _00913_ VPWR VGND sg13g2_mux2_1
X_12687_ _06479_ VPWR _06498_ VGND net1735 _06497_ sg13g2_o21ai_1
X_11707_ _05611_ _05601_ _05610_ VPWR VGND sg13g2_nand2_1
X_14426_ _00227_ VGND VPWR _00965_ fpmul.seg_reg0.q\[11\] clknet_leaf_78_clk sg13g2_dfrbpq_1
X_11638_ _05543_ _05470_ _05483_ _05506_ _05477_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_566 VPWR VGND sg13g2_decap_8
X_14357_ _00158_ VGND VPWR _00899_ _00010_ clknet_leaf_86_clk sg13g2_dfrbpq_1
X_13308_ _07018_ _06952_ _07019_ VPWR VGND sg13g2_nor2_1
XFILLER_10_290 VPWR VGND sg13g2_fill_1
X_11569_ _05474_ _05473_ _05448_ VPWR VGND sg13g2_nand2_1
XFILLER_116_649 VPWR VGND sg13g2_decap_8
XFILLER_115_126 VPWR VGND sg13g2_decap_8
X_14288_ _00089_ VGND VPWR _00001_ acc_sum.reg1en.d\[0\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_111_321 VPWR VGND sg13g2_fill_1
XFILLER_97_522 VPWR VGND sg13g2_fill_1
X_08780_ _02967_ acc_sub.add_renorm0.mantisa\[4\] _02966_ VPWR VGND sg13g2_xnor2_1
XFILLER_112_866 VPWR VGND sg13g2_decap_8
X_07800_ _02094_ _02098_ _02093_ _02099_ VPWR VGND sg13g2_nand3_1
XFILLER_97_555 VPWR VGND sg13g2_decap_8
XFILLER_111_376 VPWR VGND sg13g2_fill_1
X_07731_ _02033_ _02036_ _02037_ VPWR VGND sg13g2_nor2_1
XFILLER_65_441 VPWR VGND sg13g2_decap_4
X_07662_ _01427_ _01971_ _01972_ VPWR VGND sg13g2_nand2_1
XFILLER_25_305 VPWR VGND sg13g2_fill_1
XFILLER_25_316 VPWR VGND sg13g2_decap_8
XFILLER_111_28 VPWR VGND sg13g2_decap_8
X_07593_ _01906_ VPWR _01907_ VGND _01814_ net1686 sg13g2_o21ai_1
XFILLER_65_496 VPWR VGND sg13g2_decap_8
XFILLER_53_636 VPWR VGND sg13g2_decap_8
XFILLER_37_198 VPWR VGND sg13g2_fill_1
X_09401_ _03547_ _03425_ _03466_ VPWR VGND sg13g2_nand2b_1
XFILLER_19_880 VPWR VGND sg13g2_decap_8
XFILLER_81_978 VPWR VGND sg13g2_decap_8
XFILLER_53_669 VPWR VGND sg13g2_fill_1
X_09332_ _03483_ net1738 _03479_ _03484_ VPWR VGND sg13g2_nand3_1
XFILLER_80_499 VPWR VGND sg13g2_fill_2
XFILLER_21_500 VPWR VGND sg13g2_decap_8
X_09263_ VGND VPWR _03411_ _03413_ _03417_ _03416_ sg13g2_a21oi_1
X_09194_ _03352_ VPWR _01282_ VGND net1906 _03351_ sg13g2_o21ai_1
XFILLER_14_1000 VPWR VGND sg13g2_decap_8
X_08214_ _02467_ _02468_ _02466_ _02470_ VPWR VGND _02469_ sg13g2_nand4_1
XFILLER_119_454 VPWR VGND sg13g2_fill_2
X_08145_ _02405_ _02378_ fp16_sum_pipe.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_20_14 VPWR VGND sg13g2_decap_8
X_08076_ _02341_ _02315_ _02342_ VPWR VGND sg13g2_nor2_1
XFILLER_103_800 VPWR VGND sg13g2_fill_1
Xplace1962 net1961 net1962 VPWR VGND sg13g2_buf_2
Xplace1940 net1939 net1940 VPWR VGND sg13g2_buf_2
Xplace1951 fpmul.reg1en.d\[0\] net1951 VPWR VGND sg13g2_buf_2
XFILLER_1_927 VPWR VGND sg13g2_decap_8
XFILLER_115_693 VPWR VGND sg13g2_fill_2
XFILLER_88_533 VPWR VGND sg13g2_fill_2
XFILLER_102_332 VPWR VGND sg13g2_decap_4
X_08978_ _03164_ _03163_ _03162_ VPWR VGND sg13g2_nand2b_1
XFILLER_102_376 VPWR VGND sg13g2_fill_2
XFILLER_102_365 VPWR VGND sg13g2_decap_8
XFILLER_75_227 VPWR VGND sg13g2_decap_8
XFILLER_29_56 VPWR VGND sg13g2_decap_8
XFILLER_75_238 VPWR VGND sg13g2_fill_2
XFILLER_56_441 VPWR VGND sg13g2_decap_8
X_07929_ fp16_sum_pipe.exp_mant_logic0.b\[10\] _02203_ _02204_ VPWR VGND sg13g2_nor2_1
XFILLER_28_110 VPWR VGND sg13g2_fill_1
XFILLER_84_772 VPWR VGND sg13g2_decap_8
XFILLER_57_986 VPWR VGND sg13g2_decap_4
X_10940_ net1821 _04944_ _04942_ _04947_ VPWR VGND _04946_ sg13g2_nand4_1
XFILLER_28_154 VPWR VGND sg13g2_decap_4
XFILLER_28_165 VPWR VGND sg13g2_fill_2
XFILLER_71_455 VPWR VGND sg13g2_decap_8
XFILLER_45_77 VPWR VGND sg13g2_decap_8
X_10871_ _04883_ _04772_ fp16_res_pipe.y\[14\] VPWR VGND sg13g2_nand2_1
X_13590_ VPWR _00141_ net120 VGND sg13g2_inv_1
X_12541_ fpdiv.reg_a_out\[14\] fpdiv.reg_a_out\[13\] fpdiv.reg_a_out\[12\] fpdiv.reg_a_out\[11\]
+ _06358_ VPWR VGND sg13g2_nor4_1
XFILLER_8_504 VPWR VGND sg13g2_decap_8
XFILLER_24_393 VPWR VGND sg13g2_decap_8
X_12472_ VPWR _06313_ fpmul.seg_reg0.q\[10\] VGND sg13g2_inv_1
XFILLER_40_875 VPWR VGND sg13g2_fill_2
X_14211_ VPWR _00762_ net135 VGND sg13g2_inv_1
XFILLER_124_0 VPWR VGND sg13g2_decap_8
X_11423_ VGND VPWR _05357_ net1939 _01059_ _05358_ sg13g2_a21oi_1
XFILLER_8_559 VPWR VGND sg13g2_decap_8
XFILLER_126_925 VPWR VGND sg13g2_decap_8
XFILLER_6_49 VPWR VGND sg13g2_decap_8
XFILLER_125_457 VPWR VGND sg13g2_fill_2
X_14142_ VPWR _00693_ net134 VGND sg13g2_inv_1
X_11354_ _05307_ _05306_ net1634 VPWR VGND sg13g2_nand2_1
XFILLER_106_660 VPWR VGND sg13g2_fill_2
X_14073_ VPWR _00624_ net80 VGND sg13g2_inv_1
X_11285_ _05246_ net1635 _05245_ VPWR VGND sg13g2_nand2_1
X_10305_ _04370_ net1912 fp16_res_pipe.x2\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_4_776 VPWR VGND sg13g2_decap_8
XFILLER_4_754 VPWR VGND sg13g2_decap_8
XFILLER_3_231 VPWR VGND sg13g2_decap_8
XFILLER_112_118 VPWR VGND sg13g2_decap_8
XFILLER_106_671 VPWR VGND sg13g2_fill_1
X_13024_ _06766_ _06768_ _06791_ _06792_ VPWR VGND sg13g2_nor3_1
XFILLER_10_91 VPWR VGND sg13g2_decap_8
XFILLER_3_264 VPWR VGND sg13g2_decap_8
X_10236_ _01196_ _04307_ _04308_ VPWR VGND sg13g2_nand2_1
XFILLER_126_91 VPWR VGND sg13g2_decap_8
XFILLER_86_40 VPWR VGND sg13g2_decap_8
XFILLER_79_555 VPWR VGND sg13g2_fill_2
XFILLER_120_140 VPWR VGND sg13g2_decap_8
XFILLER_79_599 VPWR VGND sg13g2_decap_4
XFILLER_79_588 VPWR VGND sg13g2_fill_2
XFILLER_0_982 VPWR VGND sg13g2_decap_8
X_10167_ _04244_ _04246_ _04247_ VPWR VGND sg13g2_nor2_1
XFILLER_86_95 VPWR VGND sg13g2_fill_1
XFILLER_66_238 VPWR VGND sg13g2_fill_2
XFILLER_59_290 VPWR VGND sg13g2_fill_2
XFILLER_13_7 VPWR VGND sg13g2_decap_8
X_10098_ _03613_ net1703 _04182_ VPWR VGND sg13g2_nor2_1
XFILLER_47_452 VPWR VGND sg13g2_fill_1
X_13926_ VPWR _00477_ net6 VGND sg13g2_inv_1
XFILLER_19_154 VPWR VGND sg13g2_decap_8
XFILLER_74_271 VPWR VGND sg13g2_decap_8
XFILLER_63_934 VPWR VGND sg13g2_decap_8
XFILLER_62_411 VPWR VGND sg13g2_fill_1
XFILLER_62_444 VPWR VGND sg13g2_decap_4
XFILLER_16_861 VPWR VGND sg13g2_decap_8
X_13857_ VPWR _00408_ net44 VGND sg13g2_inv_1
X_12808_ _06590_ _06591_ _06580_ _00908_ VPWR VGND sg13g2_nand3_1
X_13788_ VPWR _00339_ net19 VGND sg13g2_inv_1
XFILLER_50_628 VPWR VGND sg13g2_fill_1
XFILLER_50_617 VPWR VGND sg13g2_decap_8
XFILLER_31_820 VPWR VGND sg13g2_decap_8
X_12739_ _06478_ VPWR _06541_ VGND _06507_ _06540_ sg13g2_o21ai_1
X_14409_ _00210_ VGND VPWR _00948_ fpmul.reg_a_out\[6\] clknet_leaf_95_clk sg13g2_dfrbpq_2
XFILLER_117_914 VPWR VGND sg13g2_decap_8
X_09950_ VPWR VGND _04044_ _04045_ _04043_ _03992_ _04046_ _03999_ sg13g2_a221oi_1
XFILLER_125_991 VPWR VGND sg13g2_decap_8
X_08901_ VPWR _03088_ _03010_ VGND sg13g2_inv_1
XFILLER_103_129 VPWR VGND sg13g2_decap_8
X_09881_ _03982_ VPWR _01225_ VGND net1768 _03747_ sg13g2_o21ai_1
Xclkbuf_5_12__f_clk clknet_4_6_0_clk clknet_5_12__leaf_clk VPWR VGND sg13g2_buf_8
X_08832_ _03012_ _03018_ _03008_ _03019_ VPWR VGND sg13g2_nand3_1
XFILLER_97_374 VPWR VGND sg13g2_decap_4
XFILLER_111_184 VPWR VGND sg13g2_fill_1
XFILLER_73_709 VPWR VGND sg13g2_fill_1
X_08763_ VPWR _02955_ acc_sum.exp_mant_logic0.a\[4\] VGND sg13g2_inv_1
X_07714_ _02014_ _02016_ _02020_ _02021_ VPWR VGND sg13g2_nor3_1
XFILLER_66_750 VPWR VGND sg13g2_decap_8
XFILLER_122_49 VPWR VGND sg13g2_decap_8
X_08694_ _02908_ net1668 _02767_ VPWR VGND sg13g2_nand2_1
XFILLER_65_282 VPWR VGND sg13g2_fill_1
X_07645_ _01429_ _01956_ _01957_ VPWR VGND sg13g2_nand2_1
XFILLER_54_989 VPWR VGND sg13g2_decap_4
XFILLER_15_14 VPWR VGND sg13g2_decap_8
XFILLER_26_669 VPWR VGND sg13g2_decap_8
XFILLER_90_1013 VPWR VGND sg13g2_fill_1
XFILLER_90_1002 VPWR VGND sg13g2_decap_8
X_07576_ _01834_ VPWR _01890_ VGND _01794_ _01889_ sg13g2_o21ai_1
XFILLER_41_639 VPWR VGND sg13g2_decap_8
XFILLER_40_105 VPWR VGND sg13g2_decap_8
XFILLER_34_680 VPWR VGND sg13g2_decap_8
XFILLER_25_168 VPWR VGND sg13g2_decap_8
X_09315_ _03467_ VPWR _03468_ VGND _03423_ _03421_ sg13g2_o21ai_1
X_09246_ VPWR _03400_ fp16_res_pipe.op_sign_logic0.mantisa_a\[3\] VGND sg13g2_inv_1
XFILLER_31_35 VPWR VGND sg13g2_decap_8
XFILLER_119_273 VPWR VGND sg13g2_decap_4
X_09177_ VPWR _03341_ acc_sum.exp_mant_logic0.b\[8\] VGND sg13g2_inv_1
XFILLER_108_958 VPWR VGND sg13g2_decap_8
X_08128_ _02390_ _02352_ _02389_ VPWR VGND sg13g2_nand2_1
X_08059_ _02325_ _02273_ _02324_ net1691 fp16_sum_pipe.exp_mant_logic0.a\[6\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_123_939 VPWR VGND sg13g2_decap_8
XFILLER_122_416 VPWR VGND sg13g2_decap_8
Xplace1781 net1779 net1781 VPWR VGND sg13g2_buf_1
Xplace1770 _03361_ net1770 VPWR VGND sg13g2_buf_2
XFILLER_122_449 VPWR VGND sg13g2_decap_8
Xplace1792 acc_sub.exp_mant_logic0.a\[6\] net1792 VPWR VGND sg13g2_buf_2
XFILLER_89_864 VPWR VGND sg13g2_fill_2
X_10021_ _04109_ _04010_ _04108_ VPWR VGND sg13g2_xnor2_1
XFILLER_89_886 VPWR VGND sg13g2_decap_4
XFILLER_88_385 VPWR VGND sg13g2_fill_2
XFILLER_49_739 VPWR VGND sg13g2_fill_2
XFILLER_0_267 VPWR VGND sg13g2_fill_1
XFILLER_0_278 VPWR VGND sg13g2_decap_8
XFILLER_56_21 VPWR VGND sg13g2_decap_8
X_14760_ _00561_ VGND VPWR _01284_ acc_sum.exp_mant_logic0.b\[5\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
XFILLER_29_463 VPWR VGND sg13g2_fill_1
XFILLER_91_539 VPWR VGND sg13g2_fill_2
X_13711_ VPWR _00262_ net57 VGND sg13g2_inv_1
X_11972_ fpmul.reg_b_out\[12\] fpmul.reg_a_out\[12\] _05826_ VPWR VGND sg13g2_xor2_1
XFILLER_29_474 VPWR VGND sg13g2_decap_8
XFILLER_44_466 VPWR VGND sg13g2_decap_8
X_14691_ _00492_ VGND VPWR _01219_ fp16_res_pipe.seg_reg0.q\[28\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_1
XFILLER_17_658 VPWR VGND sg13g2_decap_4
X_10923_ _04737_ VPWR _04931_ VGND _04930_ _04916_ sg13g2_o21ai_1
X_13642_ VPWR _00193_ net120 VGND sg13g2_inv_1
X_10854_ _04866_ _04748_ _04865_ VPWR VGND sg13g2_nand2_1
XFILLER_72_64 VPWR VGND sg13g2_decap_4
X_13573_ VPWR _00124_ net23 VGND sg13g2_inv_1
XFILLER_9_802 VPWR VGND sg13g2_decap_4
XFILLER_13_842 VPWR VGND sg13g2_decap_8
XFILLER_31_149 VPWR VGND sg13g2_decap_8
X_12524_ _06348_ acc_sub.x2\[5\] net1956 VPWR VGND sg13g2_nand2_1
X_10785_ _04791_ _04796_ _04797_ VPWR VGND sg13g2_nor2_1
XFILLER_8_334 VPWR VGND sg13g2_decap_8
XFILLER_9_857 VPWR VGND sg13g2_decap_8
XFILLER_12_385 VPWR VGND sg13g2_fill_2
XFILLER_12_396 VPWR VGND sg13g2_decap_8
X_12455_ _06299_ _06277_ _06298_ VPWR VGND sg13g2_xnor2_1
XFILLER_126_722 VPWR VGND sg13g2_decap_8
XFILLER_125_210 VPWR VGND sg13g2_decap_8
X_11406_ VPWR _05348_ fpdiv.div_out\[3\] VGND sg13g2_inv_1
X_12386_ VPWR _06232_ _06231_ VGND sg13g2_inv_1
XFILLER_99_617 VPWR VGND sg13g2_fill_1
X_14125_ VPWR _00676_ net117 VGND sg13g2_inv_1
X_11337_ _05288_ _05289_ _05290_ _05291_ VPWR VGND sg13g2_nor3_1
XFILLER_126_799 VPWR VGND sg13g2_decap_8
XFILLER_125_287 VPWR VGND sg13g2_decap_8
XFILLER_113_416 VPWR VGND sg13g2_fill_1
XFILLER_98_149 VPWR VGND sg13g2_decap_4
X_14056_ VPWR _00607_ net96 VGND sg13g2_inv_1
XFILLER_97_72 VPWR VGND sg13g2_fill_1
XFILLER_95_801 VPWR VGND sg13g2_decap_8
X_11268_ _05231_ _05230_ net1635 VPWR VGND sg13g2_nand2_1
XFILLER_122_994 VPWR VGND sg13g2_decap_8
XFILLER_121_471 VPWR VGND sg13g2_decap_8
X_13007_ net1853 fpmul.seg_reg0.q\[7\] _06775_ VPWR VGND sg13g2_nor2_1
X_11199_ _01091_ _05165_ _05166_ VPWR VGND sg13g2_nand2_1
XFILLER_67_525 VPWR VGND sg13g2_decap_4
X_10219_ _04293_ _04177_ net1745 VPWR VGND sg13g2_nand2_1
XFILLER_94_322 VPWR VGND sg13g2_decap_8
XFILLER_39_238 VPWR VGND sg13g2_decap_8
X_14958_ _00759_ VGND VPWR _01478_ acc_sub.add_renorm0.mantisa\[2\] clknet_5_29__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_36_934 VPWR VGND sg13g2_decap_8
XFILLER_35_422 VPWR VGND sg13g2_decap_4
X_14889_ _00690_ VGND VPWR _01409_ acc_sub.exp_mant_logic0.b\[15\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_1
X_13909_ VPWR _00460_ net16 VGND sg13g2_inv_1
X_07430_ VPWR _01763_ fpdiv.divider0.divisor\[9\] VGND sg13g2_inv_1
X_07361_ _01716_ VPWR _01472_ VGND net1798 _01715_ sg13g2_o21ai_1
XFILLER_22_149 VPWR VGND sg13g2_fill_2
X_09100_ _03282_ VPWR _01306_ VGND net1801 _03272_ sg13g2_o21ai_1
XFILLER_87_0 VPWR VGND sg13g2_decap_8
X_07292_ net1667 VPWR _01659_ VGND _01526_ _01658_ sg13g2_o21ai_1
X_09031_ VGND VPWR _03144_ net1791 _03217_ _03216_ sg13g2_a21oi_1
XFILLER_117_711 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_117_788 VPWR VGND sg13g2_decap_8
XFILLER_116_243 VPWR VGND sg13g2_decap_8
XFILLER_117_49 VPWR VGND sg13g2_decap_8
XFILLER_89_105 VPWR VGND sg13g2_decap_8
XFILLER_100_611 VPWR VGND sg13g2_decap_8
X_09864_ _03972_ net1768 acc_sum.y\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_86_834 VPWR VGND sg13g2_decap_8
X_08815_ _03002_ acc_sub.add_renorm0.mantisa\[5\] VPWR VGND sg13g2_inv_2
XFILLER_112_493 VPWR VGND sg13g2_decap_8
X_09795_ _03909_ _03907_ _03908_ VPWR VGND sg13g2_nand2_1
XFILLER_86_878 VPWR VGND sg13g2_fill_1
XFILLER_39_761 VPWR VGND sg13g2_decap_8
X_08746_ _02944_ acc\[10\] net1898 VPWR VGND sg13g2_nand2_1
X_08677_ net1816 acc_sum.add_renorm0.mantisa\[5\] _02894_ VPWR VGND sg13g2_nor2_1
XFILLER_26_35 VPWR VGND sg13g2_decap_8
XFILLER_26_433 VPWR VGND sg13g2_decap_4
XFILLER_27_967 VPWR VGND sg13g2_decap_8
X_07628_ VGND VPWR _01939_ _01941_ _01942_ _01905_ sg13g2_a21oi_1
XFILLER_41_414 VPWR VGND sg13g2_decap_8
XFILLER_14_639 VPWR VGND sg13g2_decap_8
X_07559_ VPWR _01873_ _01801_ VGND sg13g2_inv_1
XFILLER_22_650 VPWR VGND sg13g2_decap_4
XFILLER_42_56 VPWR VGND sg13g2_decap_8
X_10570_ _04598_ acc_sub.x2\[14\] net1925 VPWR VGND sg13g2_nand2_1
XFILLER_21_160 VPWR VGND sg13g2_decap_4
X_09229_ VPWR _03383_ _03382_ VGND sg13g2_inv_1
XFILLER_5_304 VPWR VGND sg13g2_fill_2
XFILLER_10_856 VPWR VGND sg13g2_decap_8
X_12240_ _06086_ _06077_ _06085_ VPWR VGND sg13g2_nand2_1
XFILLER_5_315 VPWR VGND sg13g2_fill_2
XFILLER_108_766 VPWR VGND sg13g2_fill_1
X_12171_ VPWR _06017_ _06016_ VGND sg13g2_inv_1
XFILLER_107_287 VPWR VGND sg13g2_decap_8
XFILLER_107_265 VPWR VGND sg13g2_decap_8
XFILLER_122_224 VPWR VGND sg13g2_decap_8
XFILLER_104_950 VPWR VGND sg13g2_decap_8
X_11122_ _05092_ _05009_ _05091_ acc_sum.exp_mant_logic0.b\[14\] _02935_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_95_119 VPWR VGND sg13g2_decap_8
X_11053_ VPWR _05031_ _05016_ VGND sg13g2_inv_1
XFILLER_1_587 VPWR VGND sg13g2_fill_2
XFILLER_77_834 VPWR VGND sg13g2_decap_8
XFILLER_67_64 VPWR VGND sg13g2_fill_1
XFILLER_67_53 VPWR VGND sg13g2_fill_1
X_10004_ _04092_ _03589_ fp16_res_pipe.exp_mant_logic0.b\[14\] VPWR VGND sg13g2_nand2_1
X_14812_ _00613_ VGND VPWR _01336_ acc_sum.add_renorm0.mantisa\[1\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
XFILLER_91_303 VPWR VGND sg13g2_fill_1
XFILLER_67_86 VPWR VGND sg13g2_decap_8
XFILLER_123_70 VPWR VGND sg13g2_decap_8
XFILLER_92_859 VPWR VGND sg13g2_decap_8
XFILLER_91_325 VPWR VGND sg13g2_decap_4
XFILLER_91_314 VPWR VGND sg13g2_decap_4
XFILLER_57_580 VPWR VGND sg13g2_decap_8
XFILLER_17_411 VPWR VGND sg13g2_decap_8
XFILLER_18_934 VPWR VGND sg13g2_decap_8
XFILLER_91_347 VPWR VGND sg13g2_decap_8
X_11955_ _05814_ net1882 fpmul.reg_b_out\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_33_904 VPWR VGND sg13g2_decap_8
X_14743_ _00544_ VGND VPWR _01271_ fp16_res_pipe.add_renorm0.mantisa\[6\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_2
XFILLER_83_96 VPWR VGND sg13g2_decap_8
XFILLER_45_797 VPWR VGND sg13g2_decap_8
X_14674_ _00475_ VGND VPWR _01202_ fp16_res_pipe.op_sign_logic0.mantisa_a\[0\] clknet_leaf_144_clk
+ sg13g2_dfrbpq_2
X_10906_ VPWR _04915_ _04796_ VGND sg13g2_inv_1
X_11886_ _05772_ _05773_ _01011_ VPWR VGND sg13g2_and2_1
X_13625_ VPWR _00176_ net69 VGND sg13g2_inv_1
XFILLER_60_789 VPWR VGND sg13g2_fill_2
XFILLER_34_1003 VPWR VGND sg13g2_decap_8
X_10837_ _04849_ _04802_ VPWR VGND sg13g2_inv_2
X_13556_ VPWR _00107_ net16 VGND sg13g2_inv_1
XFILLER_13_683 VPWR VGND sg13g2_decap_8
X_10768_ _03578_ _04779_ _04780_ VPWR VGND sg13g2_nor2_1
X_13487_ VPWR _00038_ net87 VGND sg13g2_inv_1
X_12507_ fpmul.reg_a_out\[12\] net1953 _06338_ VPWR VGND sg13g2_nor2_1
XFILLER_40_491 VPWR VGND sg13g2_decap_4
X_12438_ VGND VPWR _06270_ _05997_ _06284_ _06267_ sg13g2_a21oi_1
XFILLER_8_175 VPWR VGND sg13g2_decap_8
X_10699_ _04712_ _04638_ _04711_ VPWR VGND sg13g2_nand2_1
XFILLER_113_202 VPWR VGND sg13g2_decap_8
X_12369_ _06215_ net1859 net1867 VPWR VGND sg13g2_nand2_1
XFILLER_5_871 VPWR VGND sg13g2_decap_8
XFILLER_114_769 VPWR VGND sg13g2_decap_8
XFILLER_113_235 VPWR VGND sg13g2_decap_4
XFILLER_99_469 VPWR VGND sg13g2_decap_8
XFILLER_99_458 VPWR VGND sg13g2_fill_1
X_14108_ VPWR _00659_ net47 VGND sg13g2_inv_1
X_14039_ VPWR _00590_ net81 VGND sg13g2_inv_1
XFILLER_67_300 VPWR VGND sg13g2_decap_8
XFILLER_122_791 VPWR VGND sg13g2_decap_8
XFILLER_110_920 VPWR VGND sg13g2_decap_8
XFILLER_67_322 VPWR VGND sg13g2_decap_4
XFILLER_41_1007 VPWR VGND sg13g2_decap_8
XFILLER_95_664 VPWR VGND sg13g2_decap_8
X_08600_ _02822_ VPWR _02823_ VGND _02756_ _02821_ sg13g2_o21ai_1
XFILLER_110_997 VPWR VGND sg13g2_decap_8
X_09580_ _03697_ _03694_ _03696_ VPWR VGND sg13g2_nand2_1
XFILLER_95_697 VPWR VGND sg13g2_decap_8
XFILLER_83_859 VPWR VGND sg13g2_decap_8
XFILLER_82_303 VPWR VGND sg13g2_decap_8
X_08531_ VPWR _02755_ _02754_ VGND sg13g2_inv_1
XFILLER_36_764 VPWR VGND sg13g2_fill_1
XFILLER_36_753 VPWR VGND sg13g2_decap_4
XFILLER_24_904 VPWR VGND sg13g2_decap_8
X_08462_ _02677_ _02678_ _02695_ VPWR VGND sg13g2_xor2_1
XFILLER_63_572 VPWR VGND sg13g2_fill_2
XFILLER_35_274 VPWR VGND sg13g2_decap_8
X_07413_ _01750_ VPWR _01454_ VGND net1889 _01749_ sg13g2_o21ai_1
XFILLER_63_594 VPWR VGND sg13g2_decap_8
XFILLER_51_756 VPWR VGND sg13g2_decap_8
X_08393_ _02617_ VPWR _02630_ VGND _02608_ _02603_ sg13g2_o21ai_1
X_07344_ VGND VPWR _01704_ _01495_ _01705_ net1783 sg13g2_a21oi_1
XFILLER_10_119 VPWR VGND sg13g2_decap_8
XFILLER_32_992 VPWR VGND sg13g2_decap_8
X_07275_ _01643_ VPWR _01644_ VGND net1665 _01641_ sg13g2_o21ai_1
XFILLER_109_508 VPWR VGND sg13g2_decap_8
X_09014_ _03200_ _03193_ _03199_ VPWR VGND sg13g2_xnor2_1
XFILLER_117_552 VPWR VGND sg13g2_fill_2
XFILLER_3_819 VPWR VGND sg13g2_decap_8
XFILLER_104_235 VPWR VGND sg13g2_fill_1
XFILLER_104_279 VPWR VGND sg13g2_decap_4
X_09916_ fp16_res_pipe.exp_mant_logic0.a\[7\] _04012_ _04013_ VPWR VGND sg13g2_nor2_1
XFILLER_101_920 VPWR VGND sg13g2_decap_8
XFILLER_59_845 VPWR VGND sg13g2_fill_1
X_09847_ VGND VPWR _03733_ _03806_ _03957_ _03805_ sg13g2_a21oi_1
X_09778_ _03893_ _03867_ _03873_ VPWR VGND sg13g2_xnor2_1
XFILLER_101_997 VPWR VGND sg13g2_decap_8
XFILLER_74_848 VPWR VGND sg13g2_decap_8
XFILLER_73_325 VPWR VGND sg13g2_fill_1
XFILLER_73_314 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
X_08729_ _02933_ net1815 acc_sum.seg_reg0.q\[22\] VPWR VGND sg13g2_nand2_1
XFILLER_61_509 VPWR VGND sg13g2_fill_1
XFILLER_27_731 VPWR VGND sg13g2_decap_8
X_11740_ _05644_ _05642_ _05610_ VPWR VGND sg13g2_nand2_1
XFILLER_27_764 VPWR VGND sg13g2_decap_8
XFILLER_81_380 VPWR VGND sg13g2_fill_1
XFILLER_41_233 VPWR VGND sg13g2_decap_4
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_41_244 VPWR VGND sg13g2_decap_8
X_11671_ _05575_ VPWR _01028_ VGND _04389_ _05572_ sg13g2_o21ai_1
X_14390_ _00191_ VGND VPWR _00929_ div_result\[3\] clknet_leaf_84_clk sg13g2_dfrbpq_1
X_13410_ _07083_ VPWR _00798_ VGND _06980_ net1721 sg13g2_o21ai_1
XFILLER_41_299 VPWR VGND sg13g2_fill_2
XFILLER_41_288 VPWR VGND sg13g2_fill_1
XFILLER_41_277 VPWR VGND sg13g2_fill_1
X_10622_ fp16_res_pipe.add_renorm0.mantisa\[1\] _04629_ _04634_ _04635_ VPWR VGND
+ sg13g2_nor3_1
X_13341_ _07043_ VPWR _00827_ VGND _07042_ net1726 sg13g2_o21ai_1
X_10553_ _04587_ fp16_sum_pipe.add_renorm0.exp\[4\] VPWR VGND sg13g2_inv_2
XFILLER_6_635 VPWR VGND sg13g2_decap_8
XFILLER_5_112 VPWR VGND sg13g2_decap_8
XFILLER_10_675 VPWR VGND sg13g2_decap_8
XFILLER_10_686 VPWR VGND sg13g2_fill_2
X_13272_ acc\[9\] net1676 _06991_ VPWR VGND sg13g2_nor2_1
XFILLER_6_646 VPWR VGND sg13g2_fill_2
X_10484_ VPWR _04530_ _04460_ VGND sg13g2_inv_1
XFILLER_123_500 VPWR VGND sg13g2_fill_2
X_12223_ _06069_ net1860 net1863 VPWR VGND sg13g2_nand2_1
XFILLER_118_70 VPWR VGND sg13g2_decap_8
XFILLER_64_1007 VPWR VGND sg13g2_fill_2
X_12154_ _06000_ _05996_ _05998_ VPWR VGND sg13g2_nand2_1
XFILLER_123_588 VPWR VGND sg13g2_decap_8
X_11105_ _05075_ _05026_ VPWR VGND sg13g2_inv_2
XFILLER_2_863 VPWR VGND sg13g2_decap_8
XFILLER_96_439 VPWR VGND sg13g2_decap_8
X_12085_ _05931_ _05928_ _05929_ VPWR VGND sg13g2_nand2_1
XFILLER_1_373 VPWR VGND sg13g2_decap_8
XFILLER_110_249 VPWR VGND sg13g2_fill_2
XFILLER_77_675 VPWR VGND sg13g2_fill_1
XFILLER_77_664 VPWR VGND sg13g2_fill_2
X_11036_ acc_sum.exp_mant_logic0.b\[9\] _02945_ _05015_ VPWR VGND sg13g2_nor2_1
XFILLER_49_355 VPWR VGND sg13g2_decap_4
XFILLER_49_344 VPWR VGND sg13g2_fill_1
XFILLER_49_377 VPWR VGND sg13g2_fill_2
XFILLER_37_517 VPWR VGND sg13g2_decap_8
XFILLER_94_84 VPWR VGND sg13g2_decap_8
XFILLER_94_73 VPWR VGND sg13g2_fill_1
XFILLER_91_122 VPWR VGND sg13g2_decap_8
XFILLER_91_177 VPWR VGND sg13g2_decap_8
X_12987_ _06749_ _06754_ _06755_ VPWR VGND sg13g2_nor2_1
X_14726_ _00527_ VGND VPWR _01254_ fp16_res_pipe.exp_mant_logic0.a\[13\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
XFILLER_91_188 VPWR VGND sg13g2_fill_1
X_11938_ _05802_ VPWR _00988_ VGND net1874 _05801_ sg13g2_o21ai_1
XFILLER_33_745 VPWR VGND sg13g2_decap_4
X_11869_ add_result\[4\] _05481_ net1850 _01017_ VPWR VGND sg13g2_mux2_1
X_14657_ _00458_ VGND VPWR _01185_ fp16_res_pipe.exp_mant_logic0.b\[10\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
XFILLER_33_789 VPWR VGND sg13g2_fill_2
XFILLER_20_406 VPWR VGND sg13g2_decap_8
X_13608_ VPWR _00159_ net111 VGND sg13g2_inv_1
XFILLER_60_597 VPWR VGND sg13g2_decap_4
X_14588_ _00389_ VGND VPWR _01120_ fp16_sum_pipe.exp_mant_logic0.b\[15\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_1
XFILLER_20_428 VPWR VGND sg13g2_fill_1
XFILLER_119_828 VPWR VGND sg13g2_decap_8
X_13539_ VPWR _00090_ net89 VGND sg13g2_inv_1
XFILLER_13_491 VPWR VGND sg13g2_decap_8
XFILLER_64_2 VPWR VGND sg13g2_fill_1
XFILLER_127_883 VPWR VGND sg13g2_decap_8
XFILLER_5_690 VPWR VGND sg13g2_decap_4
XFILLER_101_205 VPWR VGND sg13g2_fill_2
XFILLER_99_255 VPWR VGND sg13g2_decap_4
XFILLER_59_119 VPWR VGND sg13g2_fill_2
X_09701_ VGND VPWR _03815_ net1807 _03817_ _03816_ sg13g2_a21oi_1
X_07962_ VPWR _02236_ _02198_ VGND sg13g2_inv_1
XFILLER_114_28 VPWR VGND sg13g2_decap_8
XFILLER_101_249 VPWR VGND sg13g2_fill_1
XFILLER_96_962 VPWR VGND sg13g2_decap_8
X_07893_ _02173_ VPWR _01397_ VGND net1892 _02089_ sg13g2_o21ai_1
XFILLER_56_804 VPWR VGND sg13g2_fill_1
XFILLER_110_794 VPWR VGND sg13g2_decap_8
X_09632_ _03683_ _03722_ _03741_ _03748_ _03749_ VPWR VGND sg13g2_and4_1
XFILLER_95_483 VPWR VGND sg13g2_decap_8
XFILLER_68_697 VPWR VGND sg13g2_fill_2
X_09563_ _03680_ _03679_ _03635_ VPWR VGND sg13g2_nand2_2
XFILLER_83_667 VPWR VGND sg13g2_decap_8
X_08514_ VPWR _02738_ _02737_ VGND sg13g2_inv_1
XFILLER_70_328 VPWR VGND sg13g2_decap_4
XFILLER_63_391 VPWR VGND sg13g2_decap_8
XFILLER_36_594 VPWR VGND sg13g2_fill_1
XFILLER_24_723 VPWR VGND sg13g2_decap_8
X_09494_ _03614_ acc_sub.x2\[2\] net1918 VPWR VGND sg13g2_nand2_1
X_08445_ _02679_ _02677_ _02678_ VPWR VGND sg13g2_nand2_1
XFILLER_12_918 VPWR VGND sg13g2_decap_8
X_08376_ _02617_ VPWR _02618_ VGND _02594_ _02603_ sg13g2_o21ai_1
XFILLER_51_586 VPWR VGND sg13g2_decap_4
XFILLER_23_14 VPWR VGND sg13g2_decap_8
X_07327_ _01690_ net1784 acc_sub.add_renorm0.mantisa\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_20_962 VPWR VGND sg13g2_decap_8
XFILLER_125_809 VPWR VGND sg13g2_decap_8
X_07258_ VGND VPWR _01627_ _01541_ _01628_ _01540_ sg13g2_a21oi_1
XFILLER_87_1007 VPWR VGND sg13g2_decap_8
XFILLER_124_308 VPWR VGND sg13g2_decap_8
X_07189_ acc_sub.op_sign_logic0.mantisa_a\[2\] _01560_ _01561_ VPWR VGND sg13g2_nor2_1
XFILLER_118_894 VPWR VGND sg13g2_decap_8
XFILLER_2_126 VPWR VGND sg13g2_decap_8
XFILLER_120_503 VPWR VGND sg13g2_decap_8
XFILLER_105_566 VPWR VGND sg13g2_decap_8
XFILLER_105_555 VPWR VGND sg13g2_fill_1
XFILLER_24_1002 VPWR VGND sg13g2_decap_8
XFILLER_101_750 VPWR VGND sg13g2_decap_8
XFILLER_87_951 VPWR VGND sg13g2_decap_8
XFILLER_86_450 VPWR VGND sg13g2_decap_8
XFILLER_59_664 VPWR VGND sg13g2_fill_2
XFILLER_24_1013 VPWR VGND sg13g2_fill_1
XFILLER_101_794 VPWR VGND sg13g2_decap_4
XFILLER_86_472 VPWR VGND sg13g2_fill_1
XFILLER_74_612 VPWR VGND sg13g2_fill_2
XFILLER_74_601 VPWR VGND sg13g2_fill_2
X_12910_ _06685_ net1909 fp16_res_pipe.y\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_59_697 VPWR VGND sg13g2_decap_8
XFILLER_59_675 VPWR VGND sg13g2_decap_4
XFILLER_58_174 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
X_13890_ VPWR _00441_ net49 VGND sg13g2_inv_1
X_12841_ _06622_ _06621_ net1960 VPWR VGND sg13g2_nand2_1
XFILLER_58_196 VPWR VGND sg13g2_decap_8
XFILLER_104_83 VPWR VGND sg13g2_decap_8
XFILLER_74_689 VPWR VGND sg13g2_fill_2
XFILLER_73_155 VPWR VGND sg13g2_decap_8
XFILLER_27_550 VPWR VGND sg13g2_fill_1
X_12772_ fpmul.reg3en.q\[0\] fpdiv.reg2en.q\[0\] fp16_sum_pipe.reg4en.q\[0\] load_en
+ _06557_ VPWR VGND sg13g2_nor4_1
XFILLER_64_76 VPWR VGND sg13g2_fill_2
XFILLER_54_391 VPWR VGND sg13g2_fill_2
XFILLER_54_380 VPWR VGND sg13g2_decap_8
XFILLER_42_531 VPWR VGND sg13g2_decap_8
XFILLER_14_211 VPWR VGND sg13g2_fill_2
X_14511_ _00312_ VGND VPWR _01047_ fpdiv.divider0.dividend\[6\] clknet_leaf_59_clk
+ sg13g2_dfrbpq_1
X_11723_ VGND VPWR _05626_ _05627_ _05625_ net1727 sg13g2_a21oi_2
XFILLER_15_756 VPWR VGND sg13g2_decap_8
X_14442_ _00243_ VGND VPWR _00981_ fpmul.seg_reg0.q\[27\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_9_49 VPWR VGND sg13g2_decap_8
X_11654_ _05557_ _05558_ _05556_ _05559_ VPWR VGND sg13g2_nand3_1
Xfanout92 net93 net92 VPWR VGND sg13g2_buf_1
Xfanout81 net93 net81 VPWR VGND sg13g2_buf_2
XFILLER_80_64 VPWR VGND sg13g2_decap_4
Xfanout70 net71 net70 VPWR VGND sg13g2_buf_2
X_10605_ VPWR _04618_ _04617_ VGND sg13g2_inv_1
XFILLER_80_97 VPWR VGND sg13g2_decap_8
X_14373_ _00174_ VGND VPWR _00914_ fpmul.reg_b_out\[4\] clknet_leaf_100_clk sg13g2_dfrbpq_2
XFILLER_7_944 VPWR VGND sg13g2_decap_8
XFILLER_11_973 VPWR VGND sg13g2_decap_8
X_11585_ _05449_ _05461_ _05464_ _05490_ VPWR VGND _05428_ sg13g2_nand4_1
X_13324_ VPWR _07032_ sipo.word\[14\] VGND sg13g2_inv_1
XFILLER_6_432 VPWR VGND sg13g2_decap_8
X_10536_ VGND VPWR net1670 _04500_ _04575_ net1737 sg13g2_a21oi_1
XFILLER_13_91 VPWR VGND sg13g2_decap_4
XFILLER_127_168 VPWR VGND sg13g2_decap_8
X_13255_ VPWR VGND acc_sum.y\[13\] _06977_ net1729 net1743 _06978_ sipo.word\[13\]
+ sg13g2_a221oi_1
X_10467_ _04514_ VPWR _04515_ VGND _04411_ _04513_ sg13g2_o21ai_1
X_12206_ _06052_ _06050_ _06051_ VPWR VGND sg13g2_nand2_1
XFILLER_124_886 VPWR VGND sg13g2_decap_8
X_13186_ VPWR _06925_ sipo.shift_reg\[9\] VGND sg13g2_inv_1
XFILLER_43_7 VPWR VGND sg13g2_decap_8
X_10398_ VPWR _04448_ _04447_ VGND sg13g2_inv_1
XFILLER_111_514 VPWR VGND sg13g2_decap_4
X_12137_ _05982_ _05901_ _05983_ VPWR VGND sg13g2_nor2_1
XFILLER_96_258 VPWR VGND sg13g2_decap_8
X_12068_ _05914_ _05912_ _05913_ VPWR VGND sg13g2_nand2_1
XFILLER_77_461 VPWR VGND sg13g2_decap_8
XFILLER_65_601 VPWR VGND sg13g2_fill_1
X_11019_ _04998_ _04997_ VPWR VGND sg13g2_inv_2
XFILLER_38_848 VPWR VGND sg13g2_decap_8
XFILLER_93_954 VPWR VGND sg13g2_decap_8
XFILLER_65_645 VPWR VGND sg13g2_decap_8
XFILLER_18_550 VPWR VGND sg13g2_fill_1
X_14709_ _00510_ VGND VPWR _01237_ acc_sum.y\[12\] clknet_leaf_37_clk sg13g2_dfrbpq_1
XFILLER_21_704 VPWR VGND sg13g2_decap_8
XFILLER_33_564 VPWR VGND sg13g2_decap_8
X_08230_ _02484_ net1842 _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[8\] net1777
+ VPWR VGND sg13g2_a22oi_1
XFILLER_21_759 VPWR VGND sg13g2_decap_8
XFILLER_119_636 VPWR VGND sg13g2_decap_8
X_08161_ _02420_ net1659 fp16_sum_pipe.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_20_269 VPWR VGND sg13g2_fill_2
XFILLER_109_28 VPWR VGND sg13g2_decap_8
XFILLER_118_168 VPWR VGND sg13g2_decap_8
Xclkload40 clkload40/Y clknet_leaf_17_clk VPWR VGND sg13g2_inv_2
Xclkload62 clkload62/Y clknet_leaf_106_clk VPWR VGND sg13g2_inv_2
Xclkload51 clkload51/Y clknet_leaf_98_clk VPWR VGND sg13g2_inv_2
Xclkload84 clknet_leaf_37_clk clkload84/Y VPWR VGND sg13g2_inv_4
Xclkload95 clkload95/Y clknet_leaf_85_clk VPWR VGND sg13g2_inv_2
Xclkload73 clknet_leaf_19_clk clkload73/Y VPWR VGND sg13g2_inv_4
XFILLER_47_1013 VPWR VGND sg13g2_fill_1
XFILLER_115_886 VPWR VGND sg13g2_decap_8
XFILLER_125_49 VPWR VGND sg13g2_decap_8
X_08994_ _03157_ _03179_ _03180_ VPWR VGND sg13g2_nor2_1
XFILLER_114_374 VPWR VGND sg13g2_decap_8
XFILLER_102_514 VPWR VGND sg13g2_fill_1
X_07945_ _02217_ _02219_ _02220_ VPWR VGND sg13g2_nor2_2
XFILLER_84_910 VPWR VGND sg13g2_decap_8
XFILLER_18_14 VPWR VGND sg13g2_decap_8
XFILLER_28_314 VPWR VGND sg13g2_fill_2
XFILLER_110_580 VPWR VGND sg13g2_fill_1
X_09615_ VPWR _03732_ _03715_ VGND sg13g2_inv_1
X_07876_ _02165_ net1888 acc_sub.x2\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_84_987 VPWR VGND sg13g2_decap_8
XFILLER_83_464 VPWR VGND sg13g2_decap_8
XFILLER_28_369 VPWR VGND sg13g2_decap_8
X_09546_ _03662_ _03663_ VPWR VGND sg13g2_inv_4
XFILLER_55_177 VPWR VGND sg13g2_decap_4
XFILLER_52_851 VPWR VGND sg13g2_fill_1
XFILLER_34_35 VPWR VGND sg13g2_decap_8
XFILLER_24_553 VPWR VGND sg13g2_decap_8
XFILLER_24_564 VPWR VGND sg13g2_fill_2
X_09477_ VGND VPWR _03601_ net1919 _01249_ _03602_ sg13g2_a21oi_1
X_08428_ fpdiv.divider0.remainder_reg\[4\] _01774_ _02662_ VPWR VGND sg13g2_nor2_1
XFILLER_8_719 VPWR VGND sg13g2_decap_8
XFILLER_109_113 VPWR VGND sg13g2_decap_8
X_08359_ instr\[3\] _02601_ _02602_ VPWR VGND sg13g2_nor2_1
Xclkload1 VPWR clkload1/Y clknet_5_3__leaf_clk VGND sg13g2_inv_1
XFILLER_125_606 VPWR VGND sg13g2_decap_8
XFILLER_109_135 VPWR VGND sg13g2_decap_8
XFILLER_109_124 VPWR VGND sg13g2_fill_1
X_11370_ _03349_ _05194_ _05321_ VPWR VGND sg13g2_nor2_1
XFILLER_50_56 VPWR VGND sg13g2_decap_8
XFILLER_125_628 VPWR VGND sg13g2_fill_2
XFILLER_125_617 VPWR VGND sg13g2_fill_1
XFILLER_124_105 VPWR VGND sg13g2_decap_8
X_10321_ _04378_ net1921 fp16_res_pipe.x2\[5\] VPWR VGND sg13g2_nand2_1
X_13040_ _06763_ _06807_ _06808_ VPWR VGND sg13g2_nor2_1
XFILLER_4_958 VPWR VGND sg13g2_decap_8
XFILLER_3_413 VPWR VGND sg13g2_decap_8
XFILLER_121_812 VPWR VGND sg13g2_decap_8
XFILLER_106_864 VPWR VGND sg13g2_decap_8
XFILLER_79_726 VPWR VGND sg13g2_decap_8
X_10252_ net1829 _04128_ _04195_ _04323_ VPWR VGND sg13g2_nand3_1
XFILLER_120_311 VPWR VGND sg13g2_decap_4
X_10183_ _04262_ _04261_ net1637 VPWR VGND sg13g2_nand2_1
XFILLER_66_409 VPWR VGND sg13g2_decap_8
XFILLER_121_889 VPWR VGND sg13g2_decap_8
XFILLER_120_377 VPWR VGND sg13g2_fill_2
X_13942_ VPWR _00493_ net26 VGND sg13g2_inv_1
XFILLER_75_64 VPWR VGND sg13g2_decap_8
XFILLER_75_42 VPWR VGND sg13g2_decap_4
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_35_829 VPWR VGND sg13g2_fill_2
X_13873_ VPWR _00424_ net45 VGND sg13g2_inv_1
XFILLER_90_946 VPWR VGND sg13g2_decap_8
X_12824_ VGND VPWR acc\[12\] net1908 _06606_ net1909 sg13g2_a21oi_1
XFILLER_61_147 VPWR VGND sg13g2_decap_8
X_12755_ _06544_ VPWR _00914_ VGND net1956 _06025_ sg13g2_o21ai_1
XFILLER_15_542 VPWR VGND sg13g2_decap_4
XFILLER_91_63 VPWR VGND sg13g2_decap_8
XFILLER_42_361 VPWR VGND sg13g2_decap_8
XFILLER_42_350 VPWR VGND sg13g2_fill_2
X_11706_ _05604_ _05608_ _05610_ VPWR VGND sg13g2_nor2_1
XFILLER_15_586 VPWR VGND sg13g2_decap_8
XFILLER_91_96 VPWR VGND sg13g2_fill_2
X_12686_ _06497_ _06419_ _06461_ VPWR VGND sg13g2_xnor2_1
X_14425_ _00226_ VGND VPWR _00964_ fpmul.seg_reg0.q\[10\] clknet_leaf_78_clk sg13g2_dfrbpq_1
X_11637_ _05430_ _05468_ _05542_ VPWR VGND sg13g2_nor2_1
XFILLER_30_589 VPWR VGND sg13g2_fill_1
X_14356_ _00157_ VGND VPWR _00898_ _00009_ clknet_leaf_84_clk sg13g2_dfrbpq_1
X_11568_ _05442_ _05455_ _05473_ VPWR VGND sg13g2_nor2_1
XFILLER_115_105 VPWR VGND sg13g2_decap_8
X_13307_ _07018_ sipo.word\[1\] VPWR VGND sg13g2_inv_2
XFILLER_7_774 VPWR VGND sg13g2_decap_4
X_10519_ net1848 fp16_sum_pipe.add_renorm0.mantisa\[4\] _04561_ VPWR VGND sg13g2_nor2_1
XFILLER_6_251 VPWR VGND sg13g2_fill_1
XFILLER_6_240 VPWR VGND sg13g2_decap_8
X_14287_ _00088_ VGND VPWR _00002_ load_en clknet_leaf_52_clk sg13g2_dfrbpq_2
X_11499_ _05403_ VPWR _05404_ VGND net1841 _05402_ sg13g2_o21ai_1
XFILLER_124_672 VPWR VGND sg13g2_decap_8
XFILLER_112_845 VPWR VGND sg13g2_decap_8
XFILLER_69_225 VPWR VGND sg13g2_fill_1
X_13169_ _06913_ VPWR _00869_ VGND _06911_ net1713 sg13g2_o21ai_1
XFILLER_3_980 VPWR VGND sg13g2_decap_8
XFILLER_123_182 VPWR VGND sg13g2_decap_8
XFILLER_57_409 VPWR VGND sg13g2_decap_8
X_07730_ _02036_ _02034_ _02035_ VPWR VGND sg13g2_nand2_1
XFILLER_78_781 VPWR VGND sg13g2_fill_2
XFILLER_78_770 VPWR VGND sg13g2_decap_8
XFILLER_66_932 VPWR VGND sg13g2_fill_2
XFILLER_38_612 VPWR VGND sg13g2_decap_8
XFILLER_38_601 VPWR VGND sg13g2_fill_1
XFILLER_65_420 VPWR VGND sg13g2_decap_8
XFILLER_38_656 VPWR VGND sg13g2_fill_2
XFILLER_38_645 VPWR VGND sg13g2_decap_8
X_07661_ _01972_ acc_sub.exp_mant_logic0.a\[3\] net1672 acc_sub.op_sign_logic0.mantisa_a\[6\]
+ net1780 VPWR VGND sg13g2_a22oi_1
XFILLER_38_678 VPWR VGND sg13g2_decap_8
X_07592_ _01906_ net1686 _01881_ VPWR VGND sg13g2_nand2_1
XFILLER_81_957 VPWR VGND sg13g2_decap_8
X_09400_ _03546_ net1770 fp16_res_pipe.add_renorm0.mantisa\[4\] VPWR VGND sg13g2_nand2_1
X_09331_ _03446_ _03478_ _03477_ _03483_ VPWR VGND sg13g2_nand3_1
XFILLER_80_478 VPWR VGND sg13g2_decap_8
XFILLER_34_873 VPWR VGND sg13g2_decap_8
X_09262_ VPWR _03416_ _03415_ VGND sg13g2_inv_1
XFILLER_33_383 VPWR VGND sg13g2_fill_2
XFILLER_119_422 VPWR VGND sg13g2_decap_8
X_09193_ _03352_ acc_sub.x2\[3\] net1906 VPWR VGND sg13g2_nand2_1
X_08213_ _02469_ fp16_sum_pipe.exp_mant_logic0.b\[0\] VPWR VGND sg13g2_inv_2
XFILLER_101_1004 VPWR VGND sg13g2_decap_8
X_08144_ _01377_ _02403_ _02404_ VPWR VGND sg13g2_nand2_1
XFILLER_106_138 VPWR VGND sg13g2_decap_4
XFILLER_106_127 VPWR VGND sg13g2_decap_4
Xplace1930 net1924 net1930 VPWR VGND sg13g2_buf_2
X_08075_ _02341_ _02318_ _02319_ VPWR VGND sg13g2_nand2_1
XFILLER_122_609 VPWR VGND sg13g2_decap_8
Xplace1941 fpdiv.reg1en.d\[0\] net1941 VPWR VGND sg13g2_buf_2
Xplace1952 net1951 net1952 VPWR VGND sg13g2_buf_2
XFILLER_1_906 VPWR VGND sg13g2_decap_8
XFILLER_121_119 VPWR VGND sg13g2_decap_8
XFILLER_115_672 VPWR VGND sg13g2_decap_8
XFILLER_103_834 VPWR VGND sg13g2_decap_8
XFILLER_114_193 VPWR VGND sg13g2_decap_8
XFILLER_0_449 VPWR VGND sg13g2_decap_8
XFILLER_29_35 VPWR VGND sg13g2_decap_8
X_08977_ _03087_ _03158_ _03161_ _03163_ VPWR VGND sg13g2_nand3_1
XFILLER_57_921 VPWR VGND sg13g2_fill_1
XFILLER_69_792 VPWR VGND sg13g2_decap_8
XFILLER_56_420 VPWR VGND sg13g2_fill_2
X_07928_ VPWR _02203_ fp16_sum_pipe.exp_mant_logic0.a\[10\] VGND sg13g2_inv_1
X_07859_ VGND VPWR acc_sub.exp_mant_logic0.b\[2\] _01975_ _02153_ _02152_ sg13g2_a21oi_1
XFILLER_72_913 VPWR VGND sg13g2_decap_8
XFILLER_28_133 VPWR VGND sg13g2_decap_8
XFILLER_29_667 VPWR VGND sg13g2_fill_1
XFILLER_56_497 VPWR VGND sg13g2_decap_8
XFILLER_45_56 VPWR VGND sg13g2_decap_8
X_10870_ _04882_ _04856_ _04881_ VPWR VGND sg13g2_nand2_1
XFILLER_16_317 VPWR VGND sg13g2_decap_8
X_09529_ _03633_ _03635_ _03641_ _03645_ _03646_ VPWR VGND sg13g2_nor4_1
XFILLER_43_147 VPWR VGND sg13g2_fill_2
XFILLER_43_169 VPWR VGND sg13g2_decap_8
XFILLER_40_821 VPWR VGND sg13g2_fill_1
X_12540_ fpdiv.reg_a_out\[10\] fpdiv.reg_a_out\[9\] fpdiv.reg_a_out\[8\] fpdiv.reg_a_out\[7\]
+ _06357_ VPWR VGND sg13g2_nor4_1
XFILLER_61_22 VPWR VGND sg13g2_fill_2
XFILLER_40_832 VPWR VGND sg13g2_fill_1
X_12471_ _06312_ VPWR _00965_ VGND net1871 _06304_ sg13g2_o21ai_1
XFILLER_40_887 VPWR VGND sg13g2_decap_8
X_14210_ VPWR _00761_ net135 VGND sg13g2_inv_1
XFILLER_126_904 VPWR VGND sg13g2_decap_8
X_11422_ net1939 fpdiv.reg_a_out\[14\] _05358_ VPWR VGND sg13g2_nor2_1
XFILLER_61_88 VPWR VGND sg13g2_decap_8
XFILLER_117_0 VPWR VGND sg13g2_decap_8
X_14141_ VPWR _00692_ net134 VGND sg13g2_inv_1
XFILLER_6_28 VPWR VGND sg13g2_decap_8
X_11353_ _05304_ _05305_ _05300_ _05306_ VPWR VGND sg13g2_nand3_1
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_3_210 VPWR VGND sg13g2_fill_2
XFILLER_106_650 VPWR VGND sg13g2_decap_4
X_14072_ VPWR _00623_ net94 VGND sg13g2_inv_1
X_11284_ _05243_ _05244_ _05242_ _05245_ VPWR VGND sg13g2_nand3_1
X_10304_ fp16_res_pipe.exp_mant_logic0.b\[14\] fp16_res_pipe.x2\[14\] net1913 _01189_
+ VPWR VGND sg13g2_mux2_1
XFILLER_79_534 VPWR VGND sg13g2_fill_1
X_13023_ VPWR _06791_ _06790_ VGND sg13g2_inv_1
XFILLER_10_70 VPWR VGND sg13g2_decap_8
X_10235_ _04308_ fp16_res_pipe.exp_mant_logic0.b\[2\] net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[5\]
+ _03988_ VPWR VGND sg13g2_a22oi_1
XFILLER_126_70 VPWR VGND sg13g2_decap_8
XFILLER_121_642 VPWR VGND sg13g2_decap_8
XFILLER_79_567 VPWR VGND sg13g2_decap_4
XFILLER_121_675 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_fill_1
XFILLER_0_961 VPWR VGND sg13g2_decap_8
X_10166_ _04245_ VPWR _04246_ VGND _03609_ _04227_ sg13g2_o21ai_1
XFILLER_120_196 VPWR VGND sg13g2_decap_8
X_10097_ _01208_ _04180_ _04181_ VPWR VGND sg13g2_nand2_1
X_13925_ VPWR _00476_ net7 VGND sg13g2_inv_1
XFILLER_63_924 VPWR VGND sg13g2_fill_1
XFILLER_62_423 VPWR VGND sg13g2_decap_8
X_13856_ VPWR _00407_ net44 VGND sg13g2_inv_1
X_12807_ _06591_ net1716 _00019_ VPWR VGND sg13g2_nand2_1
XFILLER_62_467 VPWR VGND sg13g2_decap_8
XFILLER_37_1001 VPWR VGND sg13g2_decap_8
XFILLER_34_147 VPWR VGND sg13g2_decap_8
XFILLER_16_840 VPWR VGND sg13g2_decap_8
X_13787_ VPWR _00338_ net74 VGND sg13g2_inv_1
XFILLER_37_1012 VPWR VGND sg13g2_fill_2
X_10999_ _04985_ VPWR _01110_ VGND net1928 _02458_ sg13g2_o21ai_1
X_12738_ _06521_ VPWR _06540_ VGND _06528_ _06458_ sg13g2_o21ai_1
XFILLER_15_394 VPWR VGND sg13g2_fill_1
X_12669_ _06484_ _06354_ div_result\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_31_865 VPWR VGND sg13g2_fill_2
X_14408_ _00209_ VGND VPWR _00947_ fpmul.reg_a_out\[5\] clknet_leaf_100_clk sg13g2_dfrbpq_2
XFILLER_30_375 VPWR VGND sg13g2_decap_4
XFILLER_30_397 VPWR VGND sg13g2_decap_8
XFILLER_116_447 VPWR VGND sg13g2_fill_2
X_14339_ _00140_ VGND VPWR _00881_ fpmul.reg_p_out\[3\] clknet_leaf_82_clk sg13g2_dfrbpq_1
XFILLER_125_970 VPWR VGND sg13g2_decap_8
XFILLER_89_309 VPWR VGND sg13g2_decap_8
X_08900_ VPWR _03087_ _03017_ VGND sg13g2_inv_1
XFILLER_103_108 VPWR VGND sg13g2_decap_8
X_09880_ _03982_ net1768 acc_sum.y\[0\] VPWR VGND sg13g2_nand2_1
X_08831_ _03018_ _03004_ _03017_ _02971_ _03014_ VPWR VGND sg13g2_a22oi_1
XFILLER_106_29 VPWR VGND sg13g2_decap_8
XFILLER_98_854 VPWR VGND sg13g2_decap_4
XFILLER_97_353 VPWR VGND sg13g2_decap_8
XFILLER_32_0 VPWR VGND sg13g2_decap_8
XFILLER_100_826 VPWR VGND sg13g2_fill_2
XFILLER_98_898 VPWR VGND sg13g2_decap_8
XFILLER_39_910 VPWR VGND sg13g2_fill_2
XFILLER_111_196 VPWR VGND sg13g2_fill_2
XFILLER_100_837 VPWR VGND sg13g2_decap_8
XFILLER_97_397 VPWR VGND sg13g2_decap_8
X_08762_ _02954_ VPWR _01316_ VGND net1905 _02953_ sg13g2_o21ai_1
XFILLER_122_28 VPWR VGND sg13g2_decap_8
X_07713_ _02020_ _02017_ _02019_ VPWR VGND sg13g2_nand2_1
X_08693_ VPWR _02907_ _02821_ VGND sg13g2_inv_1
X_07644_ _01957_ net1793 net1672 acc_sub.op_sign_logic0.mantisa_a\[8\] net1780 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_39_998 VPWR VGND sg13g2_decap_8
XFILLER_25_103 VPWR VGND sg13g2_decap_8
XFILLER_26_626 VPWR VGND sg13g2_fill_2
XFILLER_65_294 VPWR VGND sg13g2_fill_1
XFILLER_53_456 VPWR VGND sg13g2_decap_8
X_07575_ VGND VPWR _01888_ _01801_ _01889_ _01800_ sg13g2_a21oi_1
XFILLER_80_264 VPWR VGND sg13g2_fill_2
X_09314_ _03467_ _03466_ _03441_ VPWR VGND sg13g2_nand2_1
XFILLER_21_320 VPWR VGND sg13g2_fill_1
XFILLER_22_832 VPWR VGND sg13g2_fill_2
X_09245_ fp16_res_pipe.op_sign_logic0.mantisa_a\[3\] _03398_ _03399_ VPWR VGND sg13g2_nor2_1
XFILLER_33_191 VPWR VGND sg13g2_decap_8
XFILLER_21_386 VPWR VGND sg13g2_fill_1
XFILLER_22_898 VPWR VGND sg13g2_decap_8
XFILLER_31_14 VPWR VGND sg13g2_decap_8
XFILLER_119_252 VPWR VGND sg13g2_decap_8
XFILLER_108_937 VPWR VGND sg13g2_decap_8
X_09176_ _03340_ VPWR _01288_ VGND net1898 _03339_ sg13g2_o21ai_1
XFILLER_110_7 VPWR VGND sg13g2_decap_8
XFILLER_107_425 VPWR VGND sg13g2_decap_8
X_08127_ _02389_ _02384_ _02388_ VPWR VGND sg13g2_nand2_1
XFILLER_123_918 VPWR VGND sg13g2_decap_8
X_08058_ VPWR _02324_ net1652 VGND sg13g2_inv_1
Xplace1760 net1759 net1760 VPWR VGND sg13g2_buf_2
Xplace1771 _03359_ net1771 VPWR VGND sg13g2_buf_2
XFILLER_115_491 VPWR VGND sg13g2_fill_2
XFILLER_103_653 VPWR VGND sg13g2_fill_2
Xplace1793 acc_sub.exp_mant_logic0.a\[5\] net1793 VPWR VGND sg13g2_buf_2
Xplace1782 _01779_ net1782 VPWR VGND sg13g2_buf_2
XFILLER_89_843 VPWR VGND sg13g2_fill_2
XFILLER_0_246 VPWR VGND sg13g2_decap_8
XFILLER_1_769 VPWR VGND sg13g2_fill_2
XFILLER_1_758 VPWR VGND sg13g2_fill_2
X_10020_ _04107_ VPWR _04108_ VGND _04013_ net1689 sg13g2_o21ai_1
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_88_397 VPWR VGND sg13g2_decap_8
X_11971_ _05824_ _05823_ _05825_ VPWR VGND sg13g2_xor2_1
XFILLER_72_721 VPWR VGND sg13g2_decap_8
XFILLER_56_261 VPWR VGND sg13g2_fill_1
X_13710_ VPWR _00261_ net68 VGND sg13g2_inv_1
XFILLER_44_423 VPWR VGND sg13g2_fill_1
X_10922_ _04849_ _04848_ _04930_ VPWR VGND sg13g2_nor2_1
XFILLER_72_765 VPWR VGND sg13g2_fill_2
X_14690_ _00491_ VGND VPWR _01218_ fp16_res_pipe.seg_reg0.q\[27\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
XFILLER_44_434 VPWR VGND sg13g2_decap_8
XFILLER_72_43 VPWR VGND sg13g2_fill_1
X_13641_ VPWR _00192_ net120 VGND sg13g2_inv_1
XFILLER_16_158 VPWR VGND sg13g2_decap_8
X_10853_ _04863_ _04864_ _04865_ VPWR VGND sg13g2_nor2b_1
X_13572_ VPWR _00123_ net32 VGND sg13g2_inv_1
XFILLER_25_692 VPWR VGND sg13g2_fill_1
X_10784_ VGND VPWR _04795_ _04796_ _04794_ net1709 sg13g2_a21oi_2
XFILLER_72_87 VPWR VGND sg13g2_decap_8
X_12523_ VGND VPWR _06346_ net1959 _00948_ _06347_ sg13g2_a21oi_1
XFILLER_12_353 VPWR VGND sg13g2_decap_8
XFILLER_24_191 VPWR VGND sg13g2_fill_2
XFILLER_13_898 VPWR VGND sg13g2_decap_8
X_12454_ _06298_ _06297_ _06280_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_379 VPWR VGND sg13g2_fill_1
X_11405_ _05347_ VPWR _01066_ VGND _05345_ fpdiv.divider0.en_r sg13g2_o21ai_1
X_12385_ _06216_ _06213_ _06231_ VPWR VGND sg13g2_xor2_1
XFILLER_126_778 VPWR VGND sg13g2_decap_8
X_14124_ VPWR _00675_ net129 VGND sg13g2_inv_1
X_11336_ _03351_ _05173_ _05290_ VPWR VGND sg13g2_nor2_1
XFILLER_125_266 VPWR VGND sg13g2_decap_8
XFILLER_107_992 VPWR VGND sg13g2_decap_8
XFILLER_99_629 VPWR VGND sg13g2_decap_8
XFILLER_98_128 VPWR VGND sg13g2_decap_8
XFILLER_98_117 VPWR VGND sg13g2_fill_1
X_14055_ VPWR _00606_ net79 VGND sg13g2_inv_1
XFILLER_4_585 VPWR VGND sg13g2_fill_2
XFILLER_4_574 VPWR VGND sg13g2_decap_8
XFILLER_79_320 VPWR VGND sg13g2_decap_8
X_13006_ VGND VPWR _06773_ _06774_ fpmul.seg_reg0.q\[11\] net1755 sg13g2_a21oi_2
X_11267_ _05228_ _05229_ _05225_ _05230_ VPWR VGND sg13g2_nand3_1
XFILLER_122_973 VPWR VGND sg13g2_decap_8
X_11198_ _05166_ net1810 net1680 acc_sum.op_sign_logic0.mantisa_a\[7\] net1759 VPWR
+ VGND sg13g2_a22oi_1
X_10218_ _04292_ _04165_ net1829 VPWR VGND sg13g2_nand2_1
XFILLER_39_228 VPWR VGND sg13g2_fill_2
X_10149_ _04229_ VPWR _04230_ VGND _03607_ _04227_ sg13g2_o21ai_1
XFILLER_94_356 VPWR VGND sg13g2_decap_8
XFILLER_36_913 VPWR VGND sg13g2_decap_8
X_14957_ _00758_ VGND VPWR _01477_ acc_sub.add_renorm0.mantisa\[1\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
XFILLER_94_389 VPWR VGND sg13g2_decap_8
XFILLER_90_540 VPWR VGND sg13g2_fill_1
X_14888_ _00689_ VGND VPWR _01408_ acc_sub.exp_mant_logic0.b\[14\] clknet_leaf_54_clk
+ sg13g2_dfrbpq_2
XFILLER_63_765 VPWR VGND sg13g2_decap_8
X_13908_ VPWR _00459_ net16 VGND sg13g2_inv_1
XFILLER_74_1009 VPWR VGND sg13g2_decap_4
XFILLER_51_927 VPWR VGND sg13g2_fill_1
X_13839_ VPWR _00390_ net29 VGND sg13g2_inv_1
XFILLER_35_467 VPWR VGND sg13g2_decap_4
X_07360_ _01716_ net1799 acc_sub.seg_reg0.q\[26\] VPWR VGND sg13g2_nand2_1
XFILLER_62_297 VPWR VGND sg13g2_fill_2
XFILLER_16_692 VPWR VGND sg13g2_decap_8
X_07291_ _01528_ _01630_ _01658_ VPWR VGND sg13g2_nor2_1
X_09030_ net1791 acc_sub.add_renorm0.exp\[7\] _03216_ VPWR VGND sg13g2_nor2_1
XFILLER_30_172 VPWR VGND sg13g2_decap_8
XFILLER_116_222 VPWR VGND sg13g2_decap_8
XFILLER_117_767 VPWR VGND sg13g2_decap_8
XFILLER_117_28 VPWR VGND sg13g2_decap_8
X_09932_ _04029_ _04009_ _04028_ VPWR VGND sg13g2_nand2_1
XFILLER_113_984 VPWR VGND sg13g2_decap_8
X_09863_ _03971_ VPWR _01232_ VGND acc_sum.reg3en.q\[0\] _03966_ sg13g2_o21ai_1
X_08814_ _03000_ _03001_ VPWR VGND sg13g2_inv_4
XFILLER_112_472 VPWR VGND sg13g2_decap_8
X_09794_ _03908_ _03836_ VPWR VGND sg13g2_inv_2
XFILLER_86_857 VPWR VGND sg13g2_fill_1
XFILLER_85_312 VPWR VGND sg13g2_decap_4
XFILLER_58_548 VPWR VGND sg13g2_fill_2
X_08745_ VPWR _02943_ acc_sum.exp_mant_logic0.a\[10\] VGND sg13g2_inv_1
XFILLER_39_740 VPWR VGND sg13g2_decap_8
XFILLER_26_14 VPWR VGND sg13g2_decap_8
XFILLER_27_946 VPWR VGND sg13g2_decap_8
X_08676_ _02893_ _02781_ _02892_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_294 VPWR VGND sg13g2_decap_8
X_07627_ _01941_ _01940_ _01819_ VPWR VGND sg13g2_nand2_1
XFILLER_81_573 VPWR VGND sg13g2_fill_1
XFILLER_41_404 VPWR VGND sg13g2_decap_4
XFILLER_14_618 VPWR VGND sg13g2_decap_4
XFILLER_26_478 VPWR VGND sg13g2_decap_8
XFILLER_41_448 VPWR VGND sg13g2_decap_8
XFILLER_13_139 VPWR VGND sg13g2_fill_1
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_41_459 VPWR VGND sg13g2_fill_2
XFILLER_22_640 VPWR VGND sg13g2_decap_4
X_07489_ acc_sub.exp_mant_logic0.b\[8\] acc_sub.exp_mant_logic0.a\[8\] _01812_ VPWR
+ VGND sg13g2_xor2_1
XFILLER_50_993 VPWR VGND sg13g2_fill_1
XFILLER_10_835 VPWR VGND sg13g2_decap_8
X_09228_ _03379_ _03381_ _03382_ VPWR VGND sg13g2_nor2_2
XFILLER_21_194 VPWR VGND sg13g2_decap_4
XFILLER_108_745 VPWR VGND sg13g2_decap_8
X_09159_ _03329_ acc_sum.exp_mant_logic0.b\[14\] VPWR VGND sg13g2_inv_2
XFILLER_123_704 VPWR VGND sg13g2_fill_2
XFILLER_108_778 VPWR VGND sg13g2_fill_1
XFILLER_107_244 VPWR VGND sg13g2_decap_8
X_12170_ _06015_ _05935_ _06016_ VPWR VGND sg13g2_nor2_1
XFILLER_122_203 VPWR VGND sg13g2_decap_8
X_11121_ _05091_ _05090_ _05007_ VPWR VGND sg13g2_nand2b_1
XFILLER_103_450 VPWR VGND sg13g2_decap_8
X_11052_ _05029_ VPWR _05030_ VGND _05021_ _05019_ sg13g2_o21ai_1
XFILLER_103_483 VPWR VGND sg13g2_decap_8
XFILLER_88_183 VPWR VGND sg13g2_fill_2
XFILLER_67_43 VPWR VGND sg13g2_fill_2
X_10003_ VGND VPWR _04078_ _04002_ _04091_ _03999_ sg13g2_a21oi_1
X_14811_ _00612_ VGND VPWR _01335_ acc_sum.add_renorm0.mantisa\[0\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
XFILLER_18_913 VPWR VGND sg13g2_decap_8
XFILLER_29_261 VPWR VGND sg13g2_decap_4
X_11954_ VPWR _05813_ fpmul.seg_reg0.q\[28\] VGND sg13g2_inv_1
X_14742_ _00543_ VGND VPWR _01270_ fp16_res_pipe.add_renorm0.mantisa\[5\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_2
X_11885_ _02645_ VPWR _05773_ VGND _05768_ _02654_ sg13g2_o21ai_1
XFILLER_72_562 VPWR VGND sg13g2_fill_1
XFILLER_45_776 VPWR VGND sg13g2_fill_2
XFILLER_44_253 VPWR VGND sg13g2_fill_1
X_10905_ _04914_ VPWR _01133_ VGND fp16_res_pipe.reg3en.q\[0\] _04902_ sg13g2_o21ai_1
X_14673_ _00474_ VGND VPWR _01201_ fp16_res_pipe.op_sign_logic0.mantisa_b\[10\] clknet_leaf_139_clk
+ sg13g2_dfrbpq_1
X_13624_ VPWR _00175_ net65 VGND sg13g2_inv_1
X_10836_ _04846_ _04847_ _04848_ VPWR VGND sg13g2_nor2b_1
X_13555_ VPWR _00106_ net90 VGND sg13g2_inv_1
XFILLER_41_993 VPWR VGND sg13g2_decap_8
X_10767_ _04779_ _04778_ fp16_res_pipe.add_renorm0.exp\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_73_7 VPWR VGND sg13g2_decap_4
X_13486_ VPWR _00037_ net85 VGND sg13g2_inv_1
X_12506_ VPWR _06337_ acc_sub.x2\[12\] VGND sg13g2_inv_1
XFILLER_8_154 VPWR VGND sg13g2_decap_8
XFILLER_9_655 VPWR VGND sg13g2_fill_2
X_10698_ _04711_ _04710_ _04688_ _04615_ VPWR VGND sg13g2_and3_1
X_12437_ _06283_ _06279_ _06282_ VPWR VGND sg13g2_nand2_1
XFILLER_5_850 VPWR VGND sg13g2_decap_8
X_12368_ _06214_ net1857 net1869 VPWR VGND sg13g2_nand2_1
X_14107_ VPWR _00658_ net42 VGND sg13g2_inv_1
XFILLER_114_748 VPWR VGND sg13g2_decap_8
XFILLER_99_437 VPWR VGND sg13g2_decap_8
X_12299_ _06143_ _06141_ _06145_ VPWR VGND sg13g2_nor2_1
X_11319_ _05275_ _05256_ _05274_ VPWR VGND sg13g2_nand2_1
XFILLER_122_770 VPWR VGND sg13g2_decap_8
XFILLER_101_409 VPWR VGND sg13g2_decap_8
X_14038_ VPWR _00589_ net77 VGND sg13g2_inv_1
XFILLER_80_1013 VPWR VGND sg13g2_fill_1
XFILLER_121_280 VPWR VGND sg13g2_decap_4
XFILLER_95_621 VPWR VGND sg13g2_decap_4
XFILLER_110_976 VPWR VGND sg13g2_decap_8
XFILLER_55_507 VPWR VGND sg13g2_decap_8
XFILLER_103_19 VPWR VGND sg13g2_fill_2
XFILLER_94_164 VPWR VGND sg13g2_fill_2
XFILLER_83_838 VPWR VGND sg13g2_decap_8
XFILLER_82_348 VPWR VGND sg13g2_fill_1
X_08530_ _02754_ _02747_ acc_sum.op_sign_logic0.mantisa_a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_48_592 VPWR VGND sg13g2_fill_1
XFILLER_36_743 VPWR VGND sg13g2_decap_8
X_07412_ _01750_ net1894 acc\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_51_735 VPWR VGND sg13g2_decap_8
X_08392_ _02610_ _02628_ _02629_ VPWR VGND _02618_ sg13g2_nand3b_1
XFILLER_50_256 VPWR VGND sg13g2_decap_4
X_07343_ _01703_ _01582_ _01704_ VPWR VGND sg13g2_xor2_1
XFILLER_32_971 VPWR VGND sg13g2_decap_8
X_07274_ _01643_ net1665 _01642_ VPWR VGND sg13g2_nand2_1
X_09013_ _03199_ _03197_ _03198_ VPWR VGND sg13g2_nand2_1
XFILLER_12_49 VPWR VGND sg13g2_decap_8
XFILLER_117_575 VPWR VGND sg13g2_fill_2
XFILLER_120_729 VPWR VGND sg13g2_decap_8
XFILLER_120_718 VPWR VGND sg13g2_decap_8
XFILLER_59_813 VPWR VGND sg13g2_fill_2
X_09915_ _04012_ fp16_res_pipe.exp_mant_logic0.b\[7\] VPWR VGND sg13g2_inv_2
XFILLER_113_781 VPWR VGND sg13g2_decap_8
XFILLER_100_420 VPWR VGND sg13g2_decap_4
XFILLER_99_993 VPWR VGND sg13g2_decap_8
X_09846_ VPWR _03956_ acc_sum.y\[8\] VGND sg13g2_inv_1
XFILLER_101_976 VPWR VGND sg13g2_decap_8
XFILLER_86_643 VPWR VGND sg13g2_fill_2
XFILLER_58_345 VPWR VGND sg13g2_decap_8
X_09777_ net1664 _03891_ _03890_ _03892_ VPWR VGND sg13g2_nand3_1
XFILLER_86_687 VPWR VGND sg13g2_decap_8
XFILLER_74_827 VPWR VGND sg13g2_decap_8
XFILLER_46_529 VPWR VGND sg13g2_decap_4
XFILLER_39_581 VPWR VGND sg13g2_decap_8
XFILLER_39_570 VPWR VGND sg13g2_fill_1
XFILLER_37_35 VPWR VGND sg13g2_decap_8
X_08728_ VPWR _02932_ acc_sum.add_renorm0.exp\[0\] VGND sg13g2_inv_1
X_08659_ VGND VPWR _02785_ _02741_ _02878_ _02740_ sg13g2_a21oi_1
XFILLER_26_253 VPWR VGND sg13g2_decap_4
XFILLER_26_264 VPWR VGND sg13g2_decap_4
XFILLER_41_223 VPWR VGND sg13g2_decap_8
XFILLER_15_938 VPWR VGND sg13g2_decap_8
XFILLER_26_286 VPWR VGND sg13g2_decap_8
X_11670_ _05575_ _05573_ add_result\[15\] VPWR VGND sg13g2_nand2_1
X_10621_ _04634_ _04616_ _03572_ fp16_res_pipe.add_renorm0.mantisa\[3\] _04633_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_23_982 VPWR VGND sg13g2_decap_8
X_13340_ _07043_ net1726 fp16_res_pipe.x2\[9\] VPWR VGND sg13g2_nand2_1
X_10552_ _04586_ VPWR _01158_ VGND net1846 _04585_ sg13g2_o21ai_1
X_13271_ VPWR VGND acc_sum.y\[9\] _06989_ net1729 net1743 _06990_ sipo.word\[9\] sg13g2_a221oi_1
X_12222_ _05953_ _06067_ _06068_ VPWR VGND sg13g2_nor2_1
X_10483_ VGND VPWR _04528_ net1847 _01170_ _04529_ sg13g2_a21oi_1
XFILLER_5_179 VPWR VGND sg13g2_fill_2
XFILLER_5_168 VPWR VGND sg13g2_decap_8
X_12153_ _05996_ _05998_ _05990_ _05999_ VPWR VGND sg13g2_nand3_1
XFILLER_2_842 VPWR VGND sg13g2_decap_8
XFILLER_123_567 VPWR VGND sg13g2_decap_8
XFILLER_111_729 VPWR VGND sg13g2_decap_8
XFILLER_110_206 VPWR VGND sg13g2_decap_8
X_11104_ _05074_ VPWR _01094_ VGND net1813 _02795_ sg13g2_o21ai_1
X_12084_ _05928_ _05929_ _05908_ _05930_ VPWR VGND sg13g2_nand3_1
XFILLER_1_352 VPWR VGND sg13g2_decap_8
XFILLER_110_217 VPWR VGND sg13g2_fill_1
XFILLER_104_792 VPWR VGND sg13g2_decap_8
X_11035_ _05012_ _05013_ _05014_ VPWR VGND sg13g2_nor2_1
XFILLER_49_323 VPWR VGND sg13g2_decap_8
XFILLER_92_635 VPWR VGND sg13g2_fill_2
XFILLER_92_602 VPWR VGND sg13g2_decap_8
XFILLER_49_389 VPWR VGND sg13g2_decap_8
X_12986_ VPWR _06754_ _06753_ VGND sg13g2_inv_1
XFILLER_18_721 VPWR VGND sg13g2_decap_4
XFILLER_18_754 VPWR VGND sg13g2_decap_4
XFILLER_80_819 VPWR VGND sg13g2_decap_8
X_14725_ _00526_ VGND VPWR _01253_ fp16_res_pipe.exp_mant_logic0.a\[12\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
XFILLER_60_521 VPWR VGND sg13g2_decap_8
X_11937_ _05802_ net1877 fpmul.reg_b_out\[10\] VPWR VGND sg13g2_nand2_1
X_11868_ add_result\[5\] _05515_ net1850 _01018_ VPWR VGND sg13g2_mux2_1
XFILLER_33_757 VPWR VGND sg13g2_fill_1
X_14656_ _00457_ VGND VPWR _01184_ fp16_res_pipe.exp_mant_logic0.b\[9\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_2
X_13607_ VPWR _00158_ net118 VGND sg13g2_inv_1
XFILLER_60_576 VPWR VGND sg13g2_decap_8
X_11799_ VGND VPWR net1758 _05700_ _05701_ _05572_ sg13g2_a21oi_1
XFILLER_13_470 VPWR VGND sg13g2_decap_8
XFILLER_14_993 VPWR VGND sg13g2_decap_8
X_10819_ _04831_ _04829_ _04830_ VPWR VGND sg13g2_nand2_1
X_14587_ _00388_ VGND VPWR _01119_ fp16_sum_pipe.exp_mant_logic0.b\[14\] clknet_leaf_134_clk
+ sg13g2_dfrbpq_2
XFILLER_32_267 VPWR VGND sg13g2_decap_8
XFILLER_119_807 VPWR VGND sg13g2_decap_8
X_13538_ VPWR _00089_ net87 VGND sg13g2_inv_1
XFILLER_71_4 VPWR VGND sg13g2_fill_1
XFILLER_127_862 VPWR VGND sg13g2_decap_8
X_13469_ VGND VPWR _06901_ sipo.receiving _00003_ net3 sg13g2_a21oi_1
XFILLER_126_361 VPWR VGND sg13g2_fill_2
XFILLER_114_523 VPWR VGND sg13g2_decap_8
XFILLER_102_729 VPWR VGND sg13g2_fill_1
X_07961_ VPWR _02235_ _02193_ VGND sg13g2_inv_1
XFILLER_96_941 VPWR VGND sg13g2_decap_8
X_09700_ net1807 acc_sum.add_renorm0.exp\[4\] _03816_ VPWR VGND sg13g2_nor2_1
X_07892_ _02173_ net1892 acc_sub.x2\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_67_142 VPWR VGND sg13g2_fill_2
XFILLER_110_773 VPWR VGND sg13g2_decap_8
X_09631_ _03743_ _03747_ _03748_ VPWR VGND sg13g2_nor2b_1
XFILLER_83_613 VPWR VGND sg13g2_fill_2
XFILLER_83_602 VPWR VGND sg13g2_fill_2
XFILLER_68_676 VPWR VGND sg13g2_decap_4
XFILLER_56_849 VPWR VGND sg13g2_decap_8
X_09562_ VPWR _03679_ _03658_ VGND sg13g2_inv_1
XFILLER_82_123 VPWR VGND sg13g2_decap_4
X_08513_ _02735_ _02736_ _02737_ VPWR VGND sg13g2_nor2_1
XFILLER_24_713 VPWR VGND sg13g2_fill_1
XFILLER_63_370 VPWR VGND sg13g2_decap_8
XFILLER_36_573 VPWR VGND sg13g2_decap_8
X_09493_ _03613_ fp16_res_pipe.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_inv_2
X_08444_ _02678_ fpdiv.divider0.divisor_reg\[10\] fpdiv.divider0.remainder_reg\[10\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_51_565 VPWR VGND sg13g2_decap_8
XFILLER_51_543 VPWR VGND sg13g2_decap_4
XFILLER_23_234 VPWR VGND sg13g2_fill_2
X_08375_ _02594_ _02600_ _02599_ _02617_ VPWR VGND _02611_ sg13g2_nand4_1
XFILLER_17_1010 VPWR VGND sg13g2_decap_4
XFILLER_23_267 VPWR VGND sg13g2_decap_8
X_07326_ _01688_ VPWR _01689_ VGND _01559_ _01687_ sg13g2_o21ai_1
XFILLER_104_1013 VPWR VGND sg13g2_fill_1
XFILLER_20_941 VPWR VGND sg13g2_decap_8
X_07257_ VGND VPWR _01626_ _01568_ _01627_ _01557_ sg13g2_a21oi_1
X_07188_ VPWR _01560_ acc_sub.op_sign_logic0.mantisa_b\[2\] VGND sg13g2_inv_1
XFILLER_118_873 VPWR VGND sg13g2_decap_8
XFILLER_117_361 VPWR VGND sg13g2_decap_8
XFILLER_105_534 VPWR VGND sg13g2_decap_4
XFILLER_79_908 VPWR VGND sg13g2_decap_8
XFILLER_3_639 VPWR VGND sg13g2_decap_8
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_decap_8
XFILLER_87_930 VPWR VGND sg13g2_decap_8
XFILLER_58_142 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_111_1006 VPWR VGND sg13g2_decap_8
X_09829_ net1803 _03938_ _03936_ _03941_ VPWR VGND _03940_ sg13g2_nand4_1
XFILLER_47_838 VPWR VGND sg13g2_decap_4
XFILLER_47_816 VPWR VGND sg13g2_fill_1
XFILLER_19_518 VPWR VGND sg13g2_fill_1
XFILLER_100_294 VPWR VGND sg13g2_decap_4
XFILLER_73_134 VPWR VGND sg13g2_fill_2
XFILLER_73_123 VPWR VGND sg13g2_decap_4
X_12840_ VPWR _06621_ fpmul.reg_p_out\[11\] VGND sg13g2_inv_1
X_12771_ _06553_ _06554_ _06552_ _06556_ VPWR VGND _06555_ sg13g2_nand4_1
XFILLER_64_88 VPWR VGND sg13g2_decap_8
XFILLER_42_510 VPWR VGND sg13g2_decap_8
XFILLER_27_584 VPWR VGND sg13g2_fill_2
X_14510_ _00311_ VGND VPWR _01046_ fpdiv.divider0.dividend\[5\] clknet_leaf_58_clk
+ sg13g2_dfrbpq_2
X_11722_ fp16_sum_pipe.add_renorm0.exp\[6\] net1727 _05626_ VPWR VGND sg13g2_nor2_1
XFILLER_80_21 VPWR VGND sg13g2_decap_4
X_14441_ _00242_ VGND VPWR _00980_ fpmul.seg_reg0.q\[26\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_9_28 VPWR VGND sg13g2_decap_8
X_11653_ _05558_ _05475_ _05470_ VPWR VGND sg13g2_nand2_1
XFILLER_80_43 VPWR VGND sg13g2_decap_8
Xfanout82 net83 net82 VPWR VGND sg13g2_buf_2
Xfanout71 net72 net71 VPWR VGND sg13g2_buf_2
Xfanout60 net71 net60 VPWR VGND sg13g2_buf_1
X_14372_ _00173_ VGND VPWR _00913_ fpmul.reg_b_out\[3\] clknet_leaf_106_clk sg13g2_dfrbpq_1
XFILLER_11_952 VPWR VGND sg13g2_decap_8
X_10604_ _04617_ net1823 fp16_res_pipe.add_renorm0.mantisa\[4\] VPWR VGND sg13g2_nand2_1
Xfanout93 net141 net93 VPWR VGND sg13g2_buf_2
X_13323_ _07031_ VPWR _00833_ VGND _07026_ net1725 sg13g2_o21ai_1
XFILLER_7_923 VPWR VGND sg13g2_decap_8
XFILLER_10_451 VPWR VGND sg13g2_fill_2
X_11584_ _05483_ _05465_ _05488_ _05489_ VPWR VGND sg13g2_nor3_2
XFILLER_127_147 VPWR VGND sg13g2_decap_8
X_10535_ _04574_ net1673 _04414_ VPWR VGND sg13g2_nand2b_1
XFILLER_13_70 VPWR VGND sg13g2_decap_8
X_13254_ _03244_ _02576_ _06977_ VPWR VGND sg13g2_nor2_1
XFILLER_89_52 VPWR VGND sg13g2_decap_8
X_10466_ VGND VPWR _04405_ _04400_ _04514_ _04399_ sg13g2_a21oi_1
X_12205_ _06048_ _06026_ _06046_ _06051_ VPWR VGND sg13g2_nand3_1
X_13185_ _06924_ VPWR _00864_ VGND _06923_ net1715 sg13g2_o21ai_1
XFILLER_6_488 VPWR VGND sg13g2_decap_8
XFILLER_124_865 VPWR VGND sg13g2_decap_8
XFILLER_123_353 VPWR VGND sg13g2_fill_2
XFILLER_89_96 VPWR VGND sg13g2_decap_4
X_12136_ _05982_ fpmul.reg_a_out\[6\] fpmul.reg_b_out\[4\] VPWR VGND sg13g2_nand2_1
X_10397_ _04447_ _04445_ _04446_ VPWR VGND sg13g2_nand2_1
XFILLER_123_375 VPWR VGND sg13g2_decap_4
XFILLER_36_7 VPWR VGND sg13g2_decap_8
XFILLER_111_559 VPWR VGND sg13g2_decap_4
XFILLER_78_974 VPWR VGND sg13g2_decap_8
X_12067_ VPWR _05913_ fpmul.reg_a_out\[2\] VGND sg13g2_inv_1
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_93_933 VPWR VGND sg13g2_decap_8
XFILLER_78_996 VPWR VGND sg13g2_fill_2
X_11018_ _04997_ acc_sum.exp_mant_logic0.a\[14\] acc_sum.exp_mant_logic0.b\[14\] VPWR
+ VGND sg13g2_xnor2_1
XFILLER_38_816 VPWR VGND sg13g2_decap_8
XFILLER_37_348 VPWR VGND sg13g2_decap_4
XFILLER_64_167 VPWR VGND sg13g2_fill_1
X_12969_ acc\[0\] net1907 _03983_ _06739_ VPWR VGND sg13g2_nand3_1
XFILLER_18_573 VPWR VGND sg13g2_decap_8
XFILLER_18_584 VPWR VGND sg13g2_fill_1
XFILLER_127_1013 VPWR VGND sg13g2_fill_1
XFILLER_127_1002 VPWR VGND sg13g2_decap_8
X_14708_ _00509_ VGND VPWR _01236_ acc_sum.y\[11\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_33_532 VPWR VGND sg13g2_decap_8
XFILLER_61_885 VPWR VGND sg13g2_decap_8
X_14639_ _00440_ VGND VPWR _01171_ fp16_sum_pipe.add_renorm0.mantisa\[10\] clknet_leaf_110_clk
+ sg13g2_dfrbpq_1
XFILLER_20_204 VPWR VGND sg13g2_decap_4
XFILLER_119_604 VPWR VGND sg13g2_fill_1
X_08160_ _01376_ _02418_ _02419_ VPWR VGND sg13g2_nand2_1
XFILLER_20_226 VPWR VGND sg13g2_decap_8
XFILLER_20_237 VPWR VGND sg13g2_fill_2
XFILLER_119_615 VPWR VGND sg13g2_fill_1
XFILLER_118_147 VPWR VGND sg13g2_decap_8
XFILLER_9_282 VPWR VGND sg13g2_decap_4
X_08091_ _02356_ net1645 fp16_sum_pipe.exp_mant_logic0.a\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_62_0 VPWR VGND sg13g2_decap_8
Xclkload30 VPWR clkload30/Y clknet_leaf_8_clk VGND sg13g2_inv_1
Xclkload52 clknet_leaf_120_clk clkload52/Y VPWR VGND sg13g2_inv_4
Xclkload41 clkload41/Y clknet_leaf_114_clk VPWR VGND sg13g2_inv_2
Xclkload85 clkload85/Y clknet_leaf_47_clk VPWR VGND sg13g2_inv_2
Xclkload96 VPWR clkload96/Y clknet_leaf_86_clk VGND sg13g2_inv_1
Xclkload74 clkload74/Y clknet_leaf_20_clk VPWR VGND sg13g2_inv_2
Xclkload63 VPWR clkload63/Y clknet_leaf_107_clk VGND sg13g2_inv_1
XFILLER_115_865 VPWR VGND sg13g2_decap_8
XFILLER_88_716 VPWR VGND sg13g2_decap_8
XFILLER_125_28 VPWR VGND sg13g2_decap_8
X_08993_ _03179_ _03177_ _03178_ VPWR VGND sg13g2_nand2_1
XFILLER_69_930 VPWR VGND sg13g2_fill_1
XFILLER_87_237 VPWR VGND sg13g2_decap_8
XFILLER_69_963 VPWR VGND sg13g2_decap_8
X_07944_ fp16_sum_pipe.exp_mant_logic0.b\[7\] _02218_ _02219_ VPWR VGND sg13g2_nor2_2
XFILLER_29_805 VPWR VGND sg13g2_fill_2
X_07875_ _02164_ VPWR _01406_ VGND net1887 _01795_ sg13g2_o21ai_1
XFILLER_56_613 VPWR VGND sg13g2_fill_2
XFILLER_56_602 VPWR VGND sg13g2_decap_8
X_09614_ _03723_ _03730_ _03731_ VPWR VGND sg13g2_nor2_1
XFILLER_95_281 VPWR VGND sg13g2_fill_2
XFILLER_84_966 VPWR VGND sg13g2_decap_8
XFILLER_56_657 VPWR VGND sg13g2_decap_8
XFILLER_55_101 VPWR VGND sg13g2_fill_1
XFILLER_56_679 VPWR VGND sg13g2_fill_1
X_09545_ _03649_ _03661_ _03662_ VPWR VGND sg13g2_nor2_2
Xclkbuf_leaf_129_clk clknet_5_3__leaf_clk clknet_leaf_129_clk VPWR VGND sg13g2_buf_8
XFILLER_37_882 VPWR VGND sg13g2_decap_8
XFILLER_36_381 VPWR VGND sg13g2_fill_2
XFILLER_34_14 VPWR VGND sg13g2_decap_8
XFILLER_24_532 VPWR VGND sg13g2_decap_8
X_09476_ net1919 fp16_res_pipe.exp_mant_logic0.a\[8\] _03602_ VPWR VGND sg13g2_nor2_1
X_08427_ _02661_ fpdiv.divider0.divisor_reg\[5\] fpdiv.divider0.remainder_reg\[5\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_51_362 VPWR VGND sg13g2_fill_1
XFILLER_24_587 VPWR VGND sg13g2_fill_1
XFILLER_51_384 VPWR VGND sg13g2_fill_1
XFILLER_11_226 VPWR VGND sg13g2_fill_1
X_08358_ VPWR _02601_ instr\[2\] VGND sg13g2_inv_1
Xclkload2 clknet_5_5__leaf_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_11_259 VPWR VGND sg13g2_decap_8
X_07309_ _01674_ _01535_ _01673_ VPWR VGND sg13g2_xnor2_1
XFILLER_50_35 VPWR VGND sg13g2_decap_8
X_08289_ _02535_ _02536_ _02537_ VPWR VGND sg13g2_nor2b_1
X_10320_ _04377_ VPWR _01181_ VGND net1919 _04302_ sg13g2_o21ai_1
XFILLER_4_937 VPWR VGND sg13g2_decap_8
X_10251_ _04322_ fp16_res_pipe.exp_mant_logic0.b\[0\] VPWR VGND sg13g2_inv_2
XFILLER_79_705 VPWR VGND sg13g2_decap_8
XFILLER_3_469 VPWR VGND sg13g2_decap_8
XFILLER_105_386 VPWR VGND sg13g2_decap_8
X_10182_ _04258_ _04260_ _04256_ _04261_ VPWR VGND sg13g2_nand3_1
XFILLER_121_868 VPWR VGND sg13g2_decap_8
XFILLER_120_356 VPWR VGND sg13g2_fill_1
XFILLER_93_207 VPWR VGND sg13g2_fill_2
XFILLER_59_451 VPWR VGND sg13g2_fill_1
X_13941_ VPWR _00492_ net25 VGND sg13g2_inv_1
XFILLER_75_955 VPWR VGND sg13g2_decap_4
XFILLER_59_484 VPWR VGND sg13g2_decap_8
XFILLER_47_646 VPWR VGND sg13g2_decap_4
XFILLER_47_657 VPWR VGND sg13g2_fill_1
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_90_925 VPWR VGND sg13g2_decap_8
XFILLER_90_903 VPWR VGND sg13g2_fill_2
XFILLER_62_605 VPWR VGND sg13g2_fill_1
XFILLER_46_167 VPWR VGND sg13g2_fill_1
XFILLER_35_819 VPWR VGND sg13g2_decap_8
X_13872_ VPWR _00423_ net45 VGND sg13g2_inv_1
XFILLER_74_498 VPWR VGND sg13g2_fill_1
X_12823_ VGND VPWR net1935 add_result\[12\] _06605_ net1943 sg13g2_a21oi_1
XFILLER_34_318 VPWR VGND sg13g2_fill_1
XFILLER_28_882 VPWR VGND sg13g2_decap_8
X_12754_ _06544_ fp16_res_pipe.x2\[4\] net1956 VPWR VGND sg13g2_nand2_1
XFILLER_43_874 VPWR VGND sg13g2_decap_8
XFILLER_15_565 VPWR VGND sg13g2_decap_8
X_12685_ VPWR _06496_ div_result\[9\] VGND sg13g2_inv_1
XFILLER_30_535 VPWR VGND sg13g2_decap_4
X_14424_ _00225_ VGND VPWR _00963_ fpmul.seg_reg0.q\[9\] clknet_leaf_78_clk sg13g2_dfrbpq_1
XFILLER_24_91 VPWR VGND sg13g2_decap_8
X_11636_ _05540_ VPWR _05541_ VGND _05524_ _05539_ sg13g2_o21ai_1
X_14355_ _00156_ VGND VPWR _00897_ _00008_ clknet_leaf_84_clk sg13g2_dfrbpq_1
X_11567_ _05472_ _05469_ _05470_ VPWR VGND sg13g2_nand2_1
X_13306_ VGND VPWR net1677 _07016_ _00836_ _07017_ sg13g2_a21oi_1
X_14286_ _00087_ VGND VPWR _07113_ fp16_res_pipe.reg1en.d\[0\] clknet_leaf_53_clk
+ sg13g2_dfrbpq_2
XFILLER_7_753 VPWR VGND sg13g2_decap_8
X_10518_ _04560_ _04436_ _04559_ VPWR VGND sg13g2_xnor2_1
X_13237_ _06962_ _06957_ _06959_ _06961_ VPWR VGND sg13g2_and3_2
X_11498_ _05403_ net1841 fp16_sum_pipe.add_renorm0.mantisa\[6\] VPWR VGND sg13g2_nand2_1
X_10449_ _04467_ _04497_ _04498_ VPWR VGND sg13g2_nor2_1
XFILLER_123_161 VPWR VGND sg13g2_decap_8
XFILLER_112_824 VPWR VGND sg13g2_decap_8
XFILLER_69_204 VPWR VGND sg13g2_decap_8
X_13168_ _06913_ net1713 sipo.word\[14\] VPWR VGND sg13g2_nand2_1
X_13099_ net1700 _06858_ _06857_ _06859_ VPWR VGND sg13g2_nand3_1
X_12119_ _05965_ _05947_ _05964_ VPWR VGND sg13g2_nand2_1
XFILLER_111_367 VPWR VGND sg13g2_decap_8
XFILLER_66_911 VPWR VGND sg13g2_decap_8
XFILLER_120_890 VPWR VGND sg13g2_decap_8
XFILLER_93_730 VPWR VGND sg13g2_fill_2
XFILLER_38_624 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
X_07660_ _01971_ _01970_ net1641 VPWR VGND sg13g2_nand2_1
XFILLER_66_988 VPWR VGND sg13g2_decap_8
XFILLER_37_145 VPWR VGND sg13g2_decap_8
X_07591_ _01905_ _01897_ _01904_ VPWR VGND sg13g2_nand2_2
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_52_137 VPWR VGND sg13g2_decap_8
XFILLER_34_852 VPWR VGND sg13g2_decap_4
X_09330_ _01276_ _03481_ _03482_ VPWR VGND sg13g2_nand2_1
XFILLER_18_381 VPWR VGND sg13g2_decap_8
X_09261_ _03415_ _03414_ fp16_res_pipe.op_sign_logic0.mantisa_a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_33_340 VPWR VGND sg13g2_decap_8
XFILLER_33_351 VPWR VGND sg13g2_fill_1
X_08212_ _02468_ fp16_sum_pipe.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_inv_2
XFILLER_21_535 VPWR VGND sg13g2_decap_4
X_09192_ _03351_ acc_sum.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_inv_2
X_08143_ _02404_ fp16_sum_pipe.exp_mant_logic0.a\[1\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[4\]
+ net1774 VPWR VGND sg13g2_a22oi_1
XFILLER_119_456 VPWR VGND sg13g2_fill_1
X_08074_ _02340_ _02338_ VPWR VGND sg13g2_inv_2
Xplace1920 net1912 net1920 VPWR VGND sg13g2_buf_2
XFILLER_20_49 VPWR VGND sg13g2_decap_8
XFILLER_115_651 VPWR VGND sg13g2_decap_8
Xplace1942 net1941 net1942 VPWR VGND sg13g2_buf_2
Xplace1953 net1952 net1953 VPWR VGND sg13g2_buf_2
Xplace1931 net1930 net1931 VPWR VGND sg13g2_buf_2
XFILLER_115_695 VPWR VGND sg13g2_fill_1
XFILLER_114_161 VPWR VGND sg13g2_decap_8
XFILLER_88_513 VPWR VGND sg13g2_decap_8
XFILLER_0_428 VPWR VGND sg13g2_decap_8
XFILLER_88_546 VPWR VGND sg13g2_decap_8
XFILLER_29_14 VPWR VGND sg13g2_decap_8
X_08976_ VGND VPWR _03087_ _03158_ _03162_ _03161_ sg13g2_a21oi_1
XFILLER_75_207 VPWR VGND sg13g2_fill_1
XFILLER_29_613 VPWR VGND sg13g2_decap_8
X_07927_ _02202_ _02191_ _02196_ _02201_ VPWR VGND sg13g2_and3_1
X_07858_ _02152_ _02150_ _02151_ VPWR VGND sg13g2_nand2_1
XFILLER_57_966 VPWR VGND sg13g2_fill_2
X_07789_ _02087_ _01821_ _02088_ VPWR VGND sg13g2_nor2_1
XFILLER_72_947 VPWR VGND sg13g2_fill_1
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_28_167 VPWR VGND sg13g2_fill_1
X_09528_ VPWR _03645_ _03644_ VGND sg13g2_inv_1
XFILLER_43_126 VPWR VGND sg13g2_decap_8
XFILLER_52_671 VPWR VGND sg13g2_decap_8
XFILLER_25_896 VPWR VGND sg13g2_decap_8
XFILLER_101_74 VPWR VGND sg13g2_fill_1
XFILLER_101_63 VPWR VGND sg13g2_decap_8
XFILLER_80_991 VPWR VGND sg13g2_decap_8
X_09459_ _03590_ VPWR _01255_ VGND net1915 _03589_ sg13g2_o21ai_1
XFILLER_12_535 VPWR VGND sg13g2_decap_8
XFILLER_12_546 VPWR VGND sg13g2_fill_2
X_12470_ _06311_ net1870 _06310_ _06312_ VPWR VGND sg13g2_nand3_1
XFILLER_8_528 VPWR VGND sg13g2_decap_8
XFILLER_12_568 VPWR VGND sg13g2_decap_4
X_11421_ _05357_ acc_sub.x2\[14\] VPWR VGND sg13g2_inv_2
XFILLER_8_539 VPWR VGND sg13g2_fill_1
X_14140_ VPWR _00691_ net131 VGND sg13g2_inv_1
X_11352_ _05305_ acc_sum.exp_mant_logic0.b\[1\] _05161_ _05146_ acc_sum.exp_mant_logic0.b\[4\]
+ VPWR VGND sg13g2_a22oi_1
X_10303_ _04369_ VPWR _01190_ VGND net1911 _03985_ sg13g2_o21ai_1
X_14071_ VPWR _00622_ net95 VGND sg13g2_inv_1
X_11283_ _05244_ acc_sum.exp_mant_logic0.a\[1\] net1661 acc_sum.exp_mant_logic0.a\[0\]
+ _05141_ VPWR VGND sg13g2_a22oi_1
XFILLER_117_1012 VPWR VGND sg13g2_fill_2
XFILLER_106_695 VPWR VGND sg13g2_fill_2
XFILLER_106_684 VPWR VGND sg13g2_decap_8
XFILLER_106_662 VPWR VGND sg13g2_fill_1
XFILLER_79_502 VPWR VGND sg13g2_decap_8
X_13022_ _06771_ _06774_ _06788_ _06790_ VPWR VGND sg13g2_nor3_1
X_10234_ _04307_ _04306_ _04272_ VPWR VGND sg13g2_nand2_1
XFILLER_121_621 VPWR VGND sg13g2_decap_8
XFILLER_105_183 VPWR VGND sg13g2_fill_2
XFILLER_0_940 VPWR VGND sg13g2_decap_8
X_10165_ _04245_ net1642 fp16_res_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_94_527 VPWR VGND sg13g2_decap_8
XFILLER_66_207 VPWR VGND sg13g2_fill_1
XFILLER_120_175 VPWR VGND sg13g2_decap_8
XFILLER_94_538 VPWR VGND sg13g2_fill_2
X_10096_ _04181_ fp16_res_pipe.exp_mant_logic0.a\[3\] net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[6\]
+ net1764 VPWR VGND sg13g2_a22oi_1
XFILLER_59_292 VPWR VGND sg13g2_fill_1
XFILLER_48_977 VPWR VGND sg13g2_fill_2
X_13924_ VPWR _00475_ net6 VGND sg13g2_inv_1
XFILLER_19_134 VPWR VGND sg13g2_decap_8
X_13855_ VPWR _00406_ net43 VGND sg13g2_inv_1
X_12806_ _06590_ _06588_ net1732 VPWR VGND sg13g2_nand2_1
XFILLER_34_126 VPWR VGND sg13g2_decap_8
X_13786_ VPWR _00337_ net126 VGND sg13g2_inv_1
X_10998_ _04985_ fp16_res_pipe.x2\[5\] net1927 VPWR VGND sg13g2_nand2_1
XFILLER_124_1005 VPWR VGND sg13g2_decap_8
X_12737_ _06539_ div_result\[0\] VPWR VGND sg13g2_inv_2
XFILLER_15_384 VPWR VGND sg13g2_decap_4
XFILLER_16_896 VPWR VGND sg13g2_decap_8
XFILLER_30_310 VPWR VGND sg13g2_fill_2
X_12668_ VGND VPWR _06468_ _06482_ _06483_ net1735 sg13g2_a21oi_1
X_14407_ _00208_ VGND VPWR _00946_ fpmul.reg_a_out\[4\] clknet_leaf_100_clk sg13g2_dfrbpq_1
X_11619_ _05524_ _05523_ net1757 VPWR VGND sg13g2_nand2_1
XFILLER_116_404 VPWR VGND sg13g2_fill_2
X_12599_ _06414_ _06408_ _06415_ VPWR VGND sg13g2_xor2_1
XFILLER_117_949 VPWR VGND sg13g2_decap_8
XFILLER_116_437 VPWR VGND sg13g2_fill_2
X_14338_ _00139_ VGND VPWR _00880_ fpmul.reg_p_out\[2\] clknet_leaf_83_clk sg13g2_dfrbpq_1
XFILLER_98_800 VPWR VGND sg13g2_fill_1
X_14269_ _00070_ VGND VPWR _00820_ fp16_res_pipe.x2\[2\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_98_833 VPWR VGND sg13g2_decap_8
XFILLER_124_492 VPWR VGND sg13g2_decap_4
X_08830_ _02997_ _03016_ _03017_ VPWR VGND sg13g2_nor2_2
XFILLER_112_643 VPWR VGND sg13g2_fill_2
XFILLER_112_632 VPWR VGND sg13g2_fill_2
XFILLER_97_321 VPWR VGND sg13g2_decap_8
XFILLER_25_0 VPWR VGND sg13g2_decap_8
XFILLER_97_387 VPWR VGND sg13g2_fill_1
X_08761_ _02954_ acc\[5\] net1901 VPWR VGND sg13g2_nand2_1
X_07712_ _02019_ _02018_ _01869_ VPWR VGND sg13g2_nand2_1
X_08692_ VGND VPWR _02905_ net1817 _01338_ _02906_ sg13g2_a21oi_1
XFILLER_39_977 VPWR VGND sg13g2_decap_8
XFILLER_26_605 VPWR VGND sg13g2_fill_1
X_07643_ _01956_ net1641 _01955_ VPWR VGND sg13g2_nand2_1
XFILLER_65_273 VPWR VGND sg13g2_decap_8
XFILLER_53_424 VPWR VGND sg13g2_decap_8
XFILLER_81_744 VPWR VGND sg13g2_decap_4
X_07574_ VPWR _01888_ _01887_ VGND sg13g2_inv_1
XFILLER_81_777 VPWR VGND sg13g2_decap_8
X_09313_ _03465_ VPWR _03466_ VGND _03400_ _03398_ sg13g2_o21ai_1
XFILLER_22_800 VPWR VGND sg13g2_fill_1
XFILLER_15_49 VPWR VGND sg13g2_decap_8
X_09244_ VPWR _03398_ fp16_res_pipe.op_sign_logic0.mantisa_b\[3\] VGND sg13g2_inv_1
XFILLER_22_855 VPWR VGND sg13g2_decap_8
XFILLER_22_866 VPWR VGND sg13g2_fill_1
X_09175_ _03340_ acc_sub.x2\[9\] net1897 VPWR VGND sg13g2_nand2_1
XFILLER_119_231 VPWR VGND sg13g2_decap_8
XFILLER_108_916 VPWR VGND sg13g2_decap_8
X_08126_ _02385_ _02386_ _02387_ _02388_ VPWR VGND sg13g2_nor3_1
XFILLER_107_437 VPWR VGND sg13g2_fill_2
XFILLER_107_448 VPWR VGND sg13g2_fill_2
XFILLER_103_7 VPWR VGND sg13g2_fill_2
XFILLER_116_982 VPWR VGND sg13g2_decap_8
Xplace1750 net1749 net1750 VPWR VGND sg13g2_buf_1
XFILLER_89_822 VPWR VGND sg13g2_decap_8
Xplace1761 net1759 net1761 VPWR VGND sg13g2_buf_2
XFILLER_0_203 VPWR VGND sg13g2_decap_8
Xplace1772 net1771 net1772 VPWR VGND sg13g2_buf_1
Xplace1783 _01492_ net1783 VPWR VGND sg13g2_buf_2
Xplace1794 acc_sub.exp_mant_logic0.b\[6\] net1794 VPWR VGND sg13g2_buf_2
XFILLER_89_866 VPWR VGND sg13g2_fill_1
XFILLER_0_225 VPWR VGND sg13g2_decap_8
XFILLER_103_687 VPWR VGND sg13g2_decap_4
XFILLER_102_142 VPWR VGND sg13g2_fill_2
XFILLER_48_207 VPWR VGND sg13g2_decap_8
X_08959_ _03145_ _02978_ acc_sub.add_renorm0.mantisa\[10\] VPWR VGND sg13g2_nand2_2
XFILLER_76_549 VPWR VGND sg13g2_decap_8
XFILLER_5_1011 VPWR VGND sg13g2_fill_2
X_11970_ _05824_ fpmul.reg_a_out\[14\] fpmul.reg_b_out\[14\] VPWR VGND sg13g2_xnor2_1
X_10921_ VPWR _04929_ fp16_res_pipe.y\[10\] VGND sg13g2_inv_1
XFILLER_17_638 VPWR VGND sg13g2_decap_4
XFILLER_71_221 VPWR VGND sg13g2_decap_8
XFILLER_16_115 VPWR VGND sg13g2_decap_8
XFILLER_112_84 VPWR VGND sg13g2_decap_8
X_13640_ VPWR _00191_ net123 VGND sg13g2_inv_1
XFILLER_72_799 VPWR VGND sg13g2_decap_8
XFILLER_72_788 VPWR VGND sg13g2_decap_8
XFILLER_71_265 VPWR VGND sg13g2_decap_8
XFILLER_71_243 VPWR VGND sg13g2_decap_4
X_10852_ _04864_ net1824 fp16_res_pipe.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
X_13571_ VPWR _00122_ net32 VGND sg13g2_inv_1
XFILLER_52_490 VPWR VGND sg13g2_decap_8
X_10783_ fp16_res_pipe.add_renorm0.exp\[4\] net1709 _04795_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_51_clk clknet_5_19__leaf_clk clknet_leaf_51_clk VPWR VGND sg13g2_buf_8
X_12522_ net1854 net1959 _06347_ VPWR VGND sg13g2_nor2_1
XFILLER_12_332 VPWR VGND sg13g2_decap_8
XFILLER_13_877 VPWR VGND sg13g2_decap_8
XFILLER_12_387 VPWR VGND sg13g2_fill_1
X_12453_ _06297_ _06252_ _06264_ VPWR VGND sg13g2_nand2_1
X_11404_ _05347_ net1718 fpdiv.div_out\[4\] VPWR VGND sg13g2_nand2_1
X_12384_ VGND VPWR _06226_ _06228_ _06230_ _06229_ sg13g2_a21oi_1
XFILLER_126_757 VPWR VGND sg13g2_decap_8
XFILLER_125_245 VPWR VGND sg13g2_decap_8
X_14123_ VPWR _00674_ net131 VGND sg13g2_inv_1
X_11335_ _05252_ _05194_ _05289_ VPWR VGND sg13g2_nor2_1
XFILLER_21_70 VPWR VGND sg13g2_decap_8
XFILLER_107_971 VPWR VGND sg13g2_decap_8
X_14054_ VPWR _00605_ net79 VGND sg13g2_inv_1
X_11266_ _05229_ net1809 _05192_ net1810 net1653 VPWR VGND sg13g2_a22oi_1
XFILLER_122_952 VPWR VGND sg13g2_decap_8
XFILLER_79_343 VPWR VGND sg13g2_decap_8
X_13005_ VPWR _06773_ _06772_ VGND sg13g2_inv_1
X_10217_ _04291_ net1688 fp16_res_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_97_96 VPWR VGND sg13g2_decap_8
XFILLER_97_85 VPWR VGND sg13g2_decap_8
X_11197_ _05165_ net1635 _05164_ VPWR VGND sg13g2_nand2_1
XFILLER_95_858 VPWR VGND sg13g2_fill_2
XFILLER_94_335 VPWR VGND sg13g2_decap_8
X_10148_ _04229_ net1642 fp16_res_pipe.exp_mant_logic0.a\[4\] VPWR VGND sg13g2_nand2_1
X_14956_ _00757_ VGND VPWR _01476_ acc_sub.add_renorm0.mantisa\[0\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_1
XFILLER_95_869 VPWR VGND sg13g2_decap_4
X_10079_ _04140_ _04165_ VPWR VGND sg13g2_inv_4
XFILLER_94_379 VPWR VGND sg13g2_decap_4
XFILLER_63_700 VPWR VGND sg13g2_decap_8
X_13907_ VPWR _00458_ net25 VGND sg13g2_inv_1
X_14887_ _00688_ VGND VPWR _01407_ acc_sub.exp_mant_logic0.b\[13\] clknet_leaf_54_clk
+ sg13g2_dfrbpq_2
XFILLER_63_755 VPWR VGND sg13g2_fill_1
XFILLER_36_969 VPWR VGND sg13g2_decap_8
XFILLER_62_254 VPWR VGND sg13g2_fill_2
X_13838_ VPWR _00389_ net54 VGND sg13g2_inv_1
XFILLER_16_660 VPWR VGND sg13g2_fill_1
XFILLER_23_608 VPWR VGND sg13g2_fill_1
X_13769_ VPWR _00320_ net109 VGND sg13g2_inv_1
XFILLER_62_276 VPWR VGND sg13g2_decap_4
XFILLER_16_671 VPWR VGND sg13g2_fill_1
X_07290_ VGND VPWR _01574_ _01527_ _01657_ _01524_ sg13g2_a21oi_1
Xclkbuf_leaf_42_clk clknet_5_23__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
XFILLER_43_490 VPWR VGND sg13g2_decap_8
XFILLER_117_746 VPWR VGND sg13g2_decap_8
XFILLER_116_201 VPWR VGND sg13g2_decap_8
XFILLER_8_881 VPWR VGND sg13g2_decap_8
XFILLER_116_278 VPWR VGND sg13g2_fill_1
X_09931_ _04017_ _04027_ _04028_ VPWR VGND sg13g2_nor2_1
XFILLER_113_963 VPWR VGND sg13g2_decap_8
XFILLER_112_451 VPWR VGND sg13g2_decap_8
X_09862_ _03971_ _03783_ _03970_ VPWR VGND sg13g2_nand2_1
XFILLER_86_814 VPWR VGND sg13g2_decap_8
X_08813_ _02966_ VPWR _03000_ VGND acc_sub.add_renorm0.mantisa\[3\] _02986_ sg13g2_o21ai_1
X_09793_ VPWR _03907_ _03881_ VGND sg13g2_inv_1
X_08744_ _02942_ VPWR _01322_ VGND net1903 _02941_ sg13g2_o21ai_1
XFILLER_73_519 VPWR VGND sg13g2_decap_8
XFILLER_39_796 VPWR VGND sg13g2_decap_4
XFILLER_38_251 VPWR VGND sg13g2_decap_8
XFILLER_26_402 VPWR VGND sg13g2_decap_4
XFILLER_26_413 VPWR VGND sg13g2_fill_1
XFILLER_27_925 VPWR VGND sg13g2_decap_8
X_08675_ _02829_ VPWR _02892_ VGND _02890_ _02891_ sg13g2_o21ai_1
X_07626_ VPWR _01940_ _01933_ VGND sg13g2_inv_1
XFILLER_53_254 VPWR VGND sg13g2_decap_8
XFILLER_42_939 VPWR VGND sg13g2_decap_8
X_07557_ _01821_ _01871_ VPWR VGND sg13g2_inv_4
XFILLER_41_427 VPWR VGND sg13g2_decap_8
XFILLER_13_118 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_33_clk clknet_5_20__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_50_961 VPWR VGND sg13g2_fill_2
XFILLER_42_14 VPWR VGND sg13g2_decap_8
X_07488_ _01811_ _01806_ _01810_ VPWR VGND sg13g2_nand2_1
XFILLER_10_814 VPWR VGND sg13g2_decap_8
X_09227_ fp16_res_pipe.op_sign_logic0.mantisa_a\[7\] _03380_ _03381_ VPWR VGND sg13g2_nor2_1
XFILLER_108_724 VPWR VGND sg13g2_decap_8
XFILLER_107_212 VPWR VGND sg13g2_decap_4
X_09158_ VGND VPWR _03327_ net1896 _01294_ _03328_ sg13g2_a21oi_1
XFILLER_6_829 VPWR VGND sg13g2_decap_8
XFILLER_5_306 VPWR VGND sg13g2_fill_1
X_09089_ _03272_ acc_sub.y\[11\] VPWR VGND sg13g2_inv_2
X_08109_ _02372_ fp16_sum_pipe.exp_mant_logic0.a\[5\] net1659 net1691 fp16_sum_pipe.exp_mant_logic0.a\[3\]
+ VPWR VGND sg13g2_a22oi_1
X_11120_ _05038_ VPWR _05090_ VGND _05000_ _05089_ sg13g2_o21ai_1
XFILLER_1_534 VPWR VGND sg13g2_decap_8
XFILLER_122_259 VPWR VGND sg13g2_decap_8
XFILLER_107_62 VPWR VGND sg13g2_decap_8
XFILLER_104_985 VPWR VGND sg13g2_decap_8
X_11051_ _05029_ _03341_ acc_sum.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_1_545 VPWR VGND sg13g2_fill_1
X_10002_ _04090_ _04002_ _04089_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_589 VPWR VGND sg13g2_fill_1
X_14810_ _00611_ VGND VPWR _01334_ acc_sum.add_renorm0.exp\[7\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_76_379 VPWR VGND sg13g2_fill_1
XFILLER_29_240 VPWR VGND sg13g2_decap_8
XFILLER_44_210 VPWR VGND sg13g2_fill_1
X_11953_ _05812_ VPWR _00983_ VGND net1883 _05811_ sg13g2_o21ai_1
X_14741_ _00542_ VGND VPWR _01269_ fp16_res_pipe.add_renorm0.mantisa\[4\] clknet_5_0__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_17_446 VPWR VGND sg13g2_decap_8
XFILLER_18_969 VPWR VGND sg13g2_decap_8
X_11884_ _05767_ VPWR _05772_ VGND _05769_ _02654_ sg13g2_o21ai_1
XFILLER_83_87 VPWR VGND sg13g2_fill_2
XFILLER_83_65 VPWR VGND sg13g2_decap_8
XFILLER_60_703 VPWR VGND sg13g2_fill_2
X_14672_ _00473_ VGND VPWR _01200_ fp16_res_pipe.op_sign_logic0.mantisa_b\[9\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_1
XFILLER_17_479 VPWR VGND sg13g2_fill_2
X_10904_ _04897_ _04913_ _04911_ _04914_ VPWR VGND sg13g2_nand3_1
XFILLER_73_1010 VPWR VGND sg13g2_decap_4
XFILLER_72_585 VPWR VGND sg13g2_fill_2
X_13623_ VPWR _00174_ net68 VGND sg13g2_inv_1
XFILLER_33_939 VPWR VGND sg13g2_decap_8
XFILLER_16_70 VPWR VGND sg13g2_decap_4
X_10835_ _04847_ _04735_ _04808_ VPWR VGND sg13g2_nand2_1
XFILLER_32_427 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_24_clk clknet_5_17__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_13_652 VPWR VGND sg13g2_fill_2
XFILLER_25_490 VPWR VGND sg13g2_fill_2
X_13554_ VPWR _00105_ net92 VGND sg13g2_inv_1
XFILLER_9_634 VPWR VGND sg13g2_fill_1
X_10766_ _03582_ _04777_ _04778_ VPWR VGND sg13g2_nor2_1
XFILLER_121_1008 VPWR VGND sg13g2_decap_4
X_13485_ VPWR _00036_ net84 VGND sg13g2_inv_1
X_12505_ VGND VPWR _05359_ net1951 _00955_ _06336_ sg13g2_a21oi_1
XFILLER_8_133 VPWR VGND sg13g2_decap_8
X_10697_ _04709_ VPWR _04710_ VGND net1826 _03512_ sg13g2_o21ai_1
XFILLER_12_184 VPWR VGND sg13g2_fill_1
XFILLER_66_7 VPWR VGND sg13g2_fill_2
X_12436_ VGND VPWR _06277_ _06280_ _06282_ _06281_ sg13g2_a21oi_1
XFILLER_9_689 VPWR VGND sg13g2_fill_2
XFILLER_126_576 VPWR VGND sg13g2_fill_2
X_12367_ _06192_ _06165_ _06213_ VPWR VGND sg13g2_xor2_1
X_14106_ VPWR _00657_ net42 VGND sg13g2_inv_1
X_12298_ _06144_ _06141_ _06143_ VPWR VGND sg13g2_nand2_1
X_11318_ _05272_ _05273_ _05271_ _05274_ VPWR VGND sg13g2_nand3_1
XFILLER_4_372 VPWR VGND sg13g2_decap_4
XFILLER_95_600 VPWR VGND sg13g2_decap_8
X_14037_ VPWR _00588_ net73 VGND sg13g2_inv_1
X_11249_ _05213_ _05211_ _05073_ VPWR VGND sg13g2_nand2_1
XFILLER_110_955 VPWR VGND sg13g2_decap_8
XFILLER_95_655 VPWR VGND sg13g2_fill_1
XFILLER_95_644 VPWR VGND sg13g2_decap_8
XFILLER_94_143 VPWR VGND sg13g2_decap_8
XFILLER_68_869 VPWR VGND sg13g2_decap_8
XFILLER_68_858 VPWR VGND sg13g2_fill_1
X_14939_ _00740_ VGND VPWR _01459_ acc_sub.exp_mant_logic0.a\[7\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_36_722 VPWR VGND sg13g2_decap_8
XFILLER_51_703 VPWR VGND sg13g2_decap_4
X_07411_ VPWR _01749_ acc_sub.exp_mant_logic0.a\[2\] VGND sg13g2_inv_1
X_08391_ _02600_ _02611_ _02599_ _02628_ VPWR VGND _02627_ sg13g2_nand4_1
XFILLER_24_939 VPWR VGND sg13g2_decap_8
X_07342_ _01702_ VPWR _01703_ VGND _01546_ net1665 sg13g2_o21ai_1
XFILLER_92_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_5_7__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
XFILLER_50_235 VPWR VGND sg13g2_decap_8
XFILLER_32_950 VPWR VGND sg13g2_decap_8
X_07273_ VGND VPWR _01632_ _01507_ _01642_ _01506_ sg13g2_a21oi_1
X_09012_ VPWR _03198_ _03153_ VGND sg13g2_inv_1
XFILLER_12_28 VPWR VGND sg13g2_decap_8
XFILLER_117_565 VPWR VGND sg13g2_decap_4
XFILLER_105_727 VPWR VGND sg13g2_fill_1
XFILLER_104_204 VPWR VGND sg13g2_decap_8
XFILLER_105_738 VPWR VGND sg13g2_decap_4
XFILLER_113_760 VPWR VGND sg13g2_decap_8
XFILLER_99_972 VPWR VGND sg13g2_decap_8
X_09914_ VPWR _04011_ _04010_ VGND sg13g2_inv_1
XFILLER_98_493 VPWR VGND sg13g2_decap_8
X_09845_ _03955_ VPWR _01234_ VGND net1820 _03945_ sg13g2_o21ai_1
XFILLER_59_836 VPWR VGND sg13g2_decap_8
XFILLER_101_955 VPWR VGND sg13g2_decap_8
XFILLER_37_14 VPWR VGND sg13g2_decap_8
X_09776_ _03891_ _03860_ _03832_ VPWR VGND sg13g2_nand2_1
XFILLER_100_487 VPWR VGND sg13g2_decap_4
XFILLER_100_454 VPWR VGND sg13g2_decap_8
XFILLER_85_165 VPWR VGND sg13g2_decap_4
XFILLER_67_880 VPWR VGND sg13g2_decap_8
XFILLER_2_1003 VPWR VGND sg13g2_decap_8
X_08727_ _02931_ VPWR _01328_ VGND net1815 _02930_ sg13g2_o21ai_1
XFILLER_85_198 VPWR VGND sg13g2_decap_8
X_08658_ VGND VPWR _02876_ _02743_ _02877_ _02740_ sg13g2_a21oi_1
XFILLER_82_872 VPWR VGND sg13g2_decap_8
XFILLER_54_541 VPWR VGND sg13g2_decap_8
XFILLER_42_714 VPWR VGND sg13g2_decap_8
XFILLER_15_917 VPWR VGND sg13g2_decap_8
XFILLER_26_232 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
X_07609_ net1660 _01922_ _01923_ VPWR VGND sg13g2_nor2b_2
XFILLER_81_371 VPWR VGND sg13g2_decap_8
XFILLER_53_35 VPWR VGND sg13g2_decap_8
XFILLER_14_427 VPWR VGND sg13g2_decap_8
XFILLER_14_438 VPWR VGND sg13g2_fill_2
X_08589_ _02811_ _02724_ _02812_ VPWR VGND sg13g2_nor2_1
XFILLER_23_961 VPWR VGND sg13g2_decap_8
X_10620_ VPWR _04633_ fp16_res_pipe.add_renorm0.mantisa\[2\] VGND sg13g2_inv_1
X_10551_ _04586_ fp16_sum_pipe.seg_reg0.q\[27\] net1846 VPWR VGND sg13g2_nand2_1
XFILLER_127_329 VPWR VGND sg13g2_decap_8
X_13270_ _03294_ _02576_ _06989_ VPWR VGND sg13g2_nor2_1
X_10482_ net1847 fp16_sum_pipe.add_renorm0.mantisa\[9\] _04529_ VPWR VGND sg13g2_nor2_1
X_12221_ _06067_ _06063_ _06066_ VPWR VGND sg13g2_xnor2_1
XFILLER_123_502 VPWR VGND sg13g2_fill_1
XFILLER_108_576 VPWR VGND sg13g2_fill_2
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_123_546 VPWR VGND sg13g2_decap_8
XFILLER_97_909 VPWR VGND sg13g2_fill_2
XFILLER_64_1009 VPWR VGND sg13g2_fill_1
X_12152_ _05993_ _05997_ _05992_ _05998_ VPWR VGND sg13g2_nand3_1
XFILLER_2_821 VPWR VGND sg13g2_decap_8
XFILLER_111_708 VPWR VGND sg13g2_decap_8
XFILLER_96_419 VPWR VGND sg13g2_fill_2
XFILLER_78_65 VPWR VGND sg13g2_fill_1
X_11103_ acc_sum.reg1en.q\[0\] _05073_ _05042_ _05074_ VPWR VGND sg13g2_nand3_1
X_12083_ _05923_ _05926_ _05921_ _05929_ VPWR VGND sg13g2_nand3_1
XFILLER_89_460 VPWR VGND sg13g2_decap_8
X_11034_ acc_sum.exp_mant_logic0.a\[10\] _03337_ _05013_ VPWR VGND sg13g2_nor2_1
XFILLER_2_898 VPWR VGND sg13g2_decap_8
XFILLER_77_688 VPWR VGND sg13g2_decap_8
XFILLER_64_316 VPWR VGND sg13g2_decap_8
XFILLER_49_379 VPWR VGND sg13g2_fill_1
XFILLER_18_700 VPWR VGND sg13g2_decap_8
XFILLER_91_113 VPWR VGND sg13g2_fill_1
X_12985_ _05868_ _06752_ _06753_ VPWR VGND sg13g2_nor2_1
XFILLER_73_861 VPWR VGND sg13g2_decap_8
X_11936_ VPWR _05801_ fpmul.seg_reg0.q\[34\] VGND sg13g2_inv_1
X_14724_ _00525_ VGND VPWR _01252_ fp16_res_pipe.exp_mant_logic0.a\[11\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
XFILLER_73_883 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_32_213 VPWR VGND sg13g2_decap_4
X_11867_ _05762_ VPWR _01019_ VGND net1756 _05551_ sg13g2_o21ai_1
X_14655_ _00456_ VGND VPWR _01183_ fp16_res_pipe.exp_mant_logic0.b\[8\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_2
X_13606_ VPWR _00157_ net123 VGND sg13g2_inv_1
X_11798_ _05700_ _05671_ _05669_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_972 VPWR VGND sg13g2_decap_8
X_14586_ _00387_ VGND VPWR _01118_ fp16_sum_pipe.exp_mant_logic0.b\[13\] clknet_leaf_118_clk
+ sg13g2_dfrbpq_2
X_10818_ _04791_ _04817_ _04830_ VPWR VGND sg13g2_nor2_1
X_13537_ VPWR _00088_ net86 VGND sg13g2_inv_1
X_10749_ _04712_ VPWR _04762_ VGND _04710_ _04761_ sg13g2_o21ai_1
XFILLER_118_329 VPWR VGND sg13g2_decap_8
XFILLER_9_486 VPWR VGND sg13g2_fill_2
XFILLER_127_841 VPWR VGND sg13g2_decap_8
X_13468_ VGND VPWR _06902_ _02582_ _00004_ net1753 sg13g2_a21oi_1
X_13399_ _07076_ _02566_ sipo.word_ready VPWR VGND sg13g2_nand2_2
X_12419_ VPWR _06265_ _06264_ VGND sg13g2_inv_1
XFILLER_126_395 VPWR VGND sg13g2_decap_8
XFILLER_99_213 VPWR VGND sg13g2_decap_4
XFILLER_114_579 VPWR VGND sg13g2_decap_8
XFILLER_114_568 VPWR VGND sg13g2_fill_1
XFILLER_114_557 VPWR VGND sg13g2_decap_8
XFILLER_102_708 VPWR VGND sg13g2_decap_8
X_07960_ _02234_ _02233_ _02202_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_4_clk clknet_5_5__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
XFILLER_4_84 VPWR VGND sg13g2_decap_8
X_07891_ _02172_ VPWR _01398_ VGND net1892 _02073_ sg13g2_o21ai_1
XFILLER_68_666 VPWR VGND sg13g2_fill_1
X_09630_ _03746_ VPWR _03747_ VGND acc_sum.seg_reg1.q\[21\] _03745_ sg13g2_o21ai_1
XFILLER_96_997 VPWR VGND sg13g2_decap_8
X_09561_ _03667_ _03677_ _03678_ VPWR VGND sg13g2_nor2b_2
XFILLER_83_647 VPWR VGND sg13g2_decap_8
X_08512_ acc_sum.op_sign_logic0.mantisa_b\[7\] acc_sum.op_sign_logic0.mantisa_a\[7\]
+ _02736_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_552 VPWR VGND sg13g2_decap_8
XFILLER_91_691 VPWR VGND sg13g2_decap_8
X_09492_ _03612_ VPWR _01244_ VGND net1918 _03611_ sg13g2_o21ai_1
X_08443_ _02676_ VPWR _02677_ VGND fpdiv.divider0.divisor_reg\[9\] _02656_ sg13g2_o21ai_1
XFILLER_23_246 VPWR VGND sg13g2_decap_4
X_08374_ VGND VPWR _02559_ _02589_ _01361_ _02616_ sg13g2_a21oi_1
XFILLER_11_419 VPWR VGND sg13g2_decap_8
X_07325_ VGND VPWR _01687_ _01559_ _01688_ _01656_ sg13g2_a21oi_1
Xclkbuf_5_18__f_clk clknet_4_9_0_clk clknet_5_18__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_920 VPWR VGND sg13g2_decap_8
XFILLER_23_49 VPWR VGND sg13g2_decap_8
X_07256_ VGND VPWR _01625_ _01564_ _01626_ _01561_ sg13g2_a21oi_1
XFILLER_118_852 VPWR VGND sg13g2_decap_8
XFILLER_20_997 VPWR VGND sg13g2_decap_8
X_07187_ _01559_ _01558_ VPWR VGND sg13g2_inv_2
XFILLER_105_513 VPWR VGND sg13g2_decap_8
XFILLER_59_633 VPWR VGND sg13g2_decap_8
XFILLER_58_121 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
X_09828_ _03663_ VPWR _03940_ VGND _03939_ _03907_ sg13g2_o21ai_1
XFILLER_100_251 VPWR VGND sg13g2_decap_8
XFILLER_87_986 VPWR VGND sg13g2_decap_8
XFILLER_74_614 VPWR VGND sg13g2_fill_1
XFILLER_74_603 VPWR VGND sg13g2_fill_1
XFILLER_46_316 VPWR VGND sg13g2_fill_1
X_09759_ _03875_ _03865_ _03874_ VPWR VGND sg13g2_xnor2_1
XFILLER_100_273 VPWR VGND sg13g2_fill_2
XFILLER_104_96 VPWR VGND sg13g2_decap_8
XFILLER_61_308 VPWR VGND sg13g2_decap_8
XFILLER_27_563 VPWR VGND sg13g2_decap_8
X_12770_ _00012_ _00011_ _00010_ _00009_ _06555_ VPWR VGND sg13g2_nor4_1
XFILLER_64_78 VPWR VGND sg13g2_fill_1
XFILLER_55_894 VPWR VGND sg13g2_fill_2
XFILLER_14_213 VPWR VGND sg13g2_fill_1
XFILLER_27_574 VPWR VGND sg13g2_fill_1
XFILLER_70_853 VPWR VGND sg13g2_decap_4
X_11721_ _05625_ fp16_sum_pipe.add_renorm0.exp\[6\] _05579_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_246 VPWR VGND sg13g2_decap_4
XFILLER_120_84 VPWR VGND sg13g2_decap_8
XFILLER_70_897 VPWR VGND sg13g2_decap_8
X_14440_ _00241_ VGND VPWR _00979_ fpmul.seg_reg0.q\[25\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_14_257 VPWR VGND sg13g2_decap_8
XFILLER_14_279 VPWR VGND sg13g2_fill_1
X_11652_ _05557_ _05469_ _05434_ VPWR VGND sg13g2_nand2_1
Xfanout83 net86 net83 VPWR VGND sg13g2_buf_2
Xfanout72 net2 net72 VPWR VGND sg13g2_buf_2
Xfanout61 net62 net61 VPWR VGND sg13g2_buf_2
X_14371_ _00172_ VGND VPWR _00912_ fpmul.reg_b_out\[2\] clknet_leaf_104_clk sg13g2_dfrbpq_1
Xfanout50 net51 net50 VPWR VGND sg13g2_buf_2
XFILLER_42_599 VPWR VGND sg13g2_decap_4
XFILLER_11_931 VPWR VGND sg13g2_decap_8
X_10603_ VPWR _04616_ net1823 VGND sg13g2_inv_1
Xfanout94 net96 net94 VPWR VGND sg13g2_buf_2
X_13322_ _07031_ net1725 fp16_res_pipe.x2\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_7_902 VPWR VGND sg13g2_decap_8
XFILLER_10_441 VPWR VGND sg13g2_decap_4
X_11583_ _05488_ _05487_ VPWR VGND sg13g2_inv_2
XFILLER_127_126 VPWR VGND sg13g2_decap_8
X_10534_ VGND VPWR _04572_ net1849 _01163_ _04573_ sg13g2_a21oi_1
XFILLER_10_474 VPWR VGND sg13g2_decap_8
XFILLER_109_874 VPWR VGND sg13g2_fill_2
XFILLER_109_863 VPWR VGND sg13g2_decap_8
XFILLER_7_979 VPWR VGND sg13g2_decap_8
X_10465_ VGND VPWR _04512_ _04440_ _04513_ _04439_ sg13g2_a21oi_1
XFILLER_6_467 VPWR VGND sg13g2_decap_8
XFILLER_124_844 VPWR VGND sg13g2_decap_8
XFILLER_89_75 VPWR VGND sg13g2_decap_8
X_12204_ _06050_ _06049_ _06026_ VPWR VGND sg13g2_nand2b_1
X_13184_ _06924_ net1715 sipo.word\[9\] VPWR VGND sg13g2_nand2_1
X_10396_ VGND VPWR _04442_ _04433_ _04446_ _04441_ sg13g2_a21oi_1
XFILLER_123_332 VPWR VGND sg13g2_decap_8
X_12135_ VPWR _05981_ _05980_ VGND sg13g2_inv_1
XFILLER_111_538 VPWR VGND sg13g2_decap_8
XFILLER_2_684 VPWR VGND sg13g2_decap_4
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_96_249 VPWR VGND sg13g2_decap_4
XFILLER_78_942 VPWR VGND sg13g2_decap_8
X_12066_ _05912_ fpmul.reg_a_out\[3\] fpmul.reg_b_out\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_29_7 VPWR VGND sg13g2_decap_8
XFILLER_93_912 VPWR VGND sg13g2_decap_8
XFILLER_65_614 VPWR VGND sg13g2_decap_8
X_11017_ acc_sum.exp_mant_logic0.b\[14\] _04993_ _04996_ VPWR VGND sg13g2_nor2_1
XFILLER_92_411 VPWR VGND sg13g2_decap_8
XFILLER_93_989 VPWR VGND sg13g2_decap_8
XFILLER_92_455 VPWR VGND sg13g2_decap_4
XFILLER_80_606 VPWR VGND sg13g2_fill_2
XFILLER_65_669 VPWR VGND sg13g2_decap_8
XFILLER_46_861 VPWR VGND sg13g2_decap_8
XFILLER_46_850 VPWR VGND sg13g2_fill_1
XFILLER_18_530 VPWR VGND sg13g2_decap_8
XFILLER_73_680 VPWR VGND sg13g2_fill_2
X_12968_ VGND VPWR net1936 add_result\[0\] _06738_ net1950 sg13g2_a21oi_1
XFILLER_46_872 VPWR VGND sg13g2_fill_1
XFILLER_33_511 VPWR VGND sg13g2_fill_1
XFILLER_33_522 VPWR VGND sg13g2_decap_4
X_14707_ _00508_ VGND VPWR _01235_ acc_sum.y\[10\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_73_691 VPWR VGND sg13g2_decap_4
X_12899_ _06674_ _06673_ fp16_sum_pipe.reg1en.d\[0\] _06675_ VPWR VGND sg13g2_a21o_2
XFILLER_60_330 VPWR VGND sg13g2_fill_1
X_11919_ _05790_ net1882 fpmul.reg_a_out\[1\] VPWR VGND sg13g2_nand2_1
X_14638_ _00439_ VGND VPWR _01170_ fp16_sum_pipe.add_renorm0.mantisa\[9\] clknet_leaf_110_clk
+ sg13g2_dfrbpq_2
XFILLER_21_739 VPWR VGND sg13g2_fill_1
X_14569_ _00370_ VGND VPWR fp16_sum_pipe.reg3en.q\[0\] fp16_sum_pipe.reg4en.q\[0\]
+ clknet_leaf_96_clk sg13g2_dfrbpq_2
XFILLER_118_126 VPWR VGND sg13g2_decap_8
X_08090_ _01382_ _02354_ _02355_ VPWR VGND sg13g2_nand2_1
Xclkload20 clknet_leaf_1_clk clkload20/Y VPWR VGND sg13g2_inv_4
Xclkload53 clknet_leaf_92_clk clkload53/X VPWR VGND sg13g2_buf_8
Xclkload31 clkload31/Y clknet_leaf_9_clk VPWR VGND sg13g2_inv_2
Xclkload42 clknet_leaf_116_clk clkload42/Y VPWR VGND sg13g2_inv_4
XFILLER_127_693 VPWR VGND sg13g2_decap_4
XFILLER_115_844 VPWR VGND sg13g2_decap_8
Xclkload86 VPWR clkload86/Y clknet_leaf_49_clk VGND sg13g2_inv_1
Xclkload75 VPWR clkload75/Y clknet_leaf_21_clk VGND sg13g2_inv_1
XFILLER_55_0 VPWR VGND sg13g2_decap_8
Xclkload64 clkload64/Y clknet_leaf_100_clk VPWR VGND sg13g2_inv_2
XFILLER_47_1004 VPWR VGND sg13g2_decap_8
XFILLER_6_990 VPWR VGND sg13g2_decap_8
XFILLER_114_343 VPWR VGND sg13g2_fill_2
Xclkload97 clknet_leaf_78_clk clkload97/X VPWR VGND sg13g2_buf_1
X_08992_ _03178_ _03086_ _03173_ VPWR VGND sg13g2_nand2_1
XFILLER_102_505 VPWR VGND sg13g2_decap_8
XFILLER_87_216 VPWR VGND sg13g2_decap_8
X_07943_ _02218_ fp16_sum_pipe.exp_mant_logic0.a\[7\] VPWR VGND sg13g2_inv_2
X_07874_ _02164_ net1888 acc_sub.x2\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_68_463 VPWR VGND sg13g2_fill_1
X_09613_ VPWR _03730_ _03729_ VGND sg13g2_inv_1
XFILLER_84_945 VPWR VGND sg13g2_decap_8
XFILLER_83_411 VPWR VGND sg13g2_decap_8
XFILLER_56_636 VPWR VGND sg13g2_decap_8
XFILLER_18_49 VPWR VGND sg13g2_decap_8
XFILLER_28_316 VPWR VGND sg13g2_fill_1
XFILLER_28_327 VPWR VGND sg13g2_decap_8
XFILLER_28_338 VPWR VGND sg13g2_fill_1
XFILLER_83_455 VPWR VGND sg13g2_decap_4
XFILLER_37_850 VPWR VGND sg13g2_fill_1
XFILLER_28_349 VPWR VGND sg13g2_fill_2
X_09544_ _03657_ _03660_ _03661_ VPWR VGND sg13g2_nor2_2
XFILLER_36_360 VPWR VGND sg13g2_decap_8
XFILLER_52_864 VPWR VGND sg13g2_decap_8
X_09475_ acc_sub.x2\[8\] _03601_ VPWR VGND sg13g2_inv_4
X_08426_ VPWR _02660_ _02659_ VGND sg13g2_inv_1
XFILLER_51_374 VPWR VGND sg13g2_decap_4
XFILLER_11_205 VPWR VGND sg13g2_decap_8
XFILLER_12_728 VPWR VGND sg13g2_decap_4
XFILLER_11_238 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_decap_8
X_08357_ instr\[7\] instr\[6\] instr\[5\] _02600_ VGND VPWR instr\[4\] sg13g2_nor4_2
Xclkload3 clknet_5_7__leaf_clk clkload3/X VPWR VGND sg13g2_buf_8
XFILLER_50_14 VPWR VGND sg13g2_decap_8
XFILLER_20_750 VPWR VGND sg13g2_fill_1
X_07308_ VGND VPWR _01628_ net1667 _01673_ _01672_ sg13g2_a21oi_1
X_08288_ _02536_ net1657 fp16_sum_pipe.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_nand2_1
X_07239_ _01610_ _01609_ _01522_ VPWR VGND sg13g2_nand2_1
XFILLER_109_159 VPWR VGND sg13g2_fill_1
XFILLER_4_916 VPWR VGND sg13g2_decap_8
X_10250_ _04320_ VPWR _04321_ VGND _04300_ _04175_ sg13g2_o21ai_1
XFILLER_59_23 VPWR VGND sg13g2_fill_1
XFILLER_3_448 VPWR VGND sg13g2_decap_8
XFILLER_59_67 VPWR VGND sg13g2_fill_2
XFILLER_59_56 VPWR VGND sg13g2_decap_8
X_10181_ VGND VPWR fp16_res_pipe.exp_mant_logic0.a\[1\] _04177_ _04260_ _04259_ sg13g2_a21oi_1
XFILLER_121_847 VPWR VGND sg13g2_decap_8
XFILLER_120_379 VPWR VGND sg13g2_fill_1
XFILLER_59_463 VPWR VGND sg13g2_decap_8
X_13940_ VPWR _00491_ net16 VGND sg13g2_inv_1
XFILLER_115_84 VPWR VGND sg13g2_decap_8
XFILLER_86_260 VPWR VGND sg13g2_fill_1
XFILLER_75_934 VPWR VGND sg13g2_fill_2
XFILLER_74_422 VPWR VGND sg13g2_decap_4
XFILLER_47_625 VPWR VGND sg13g2_decap_8
XFILLER_19_327 VPWR VGND sg13g2_decap_8
X_13871_ VPWR _00422_ net45 VGND sg13g2_inv_1
XFILLER_28_850 VPWR VGND sg13g2_fill_1
X_12822_ _00018_ net1730 net1701 _06604_ VPWR VGND sg13g2_nand3_1
XFILLER_74_477 VPWR VGND sg13g2_decap_4
XFILLER_62_639 VPWR VGND sg13g2_decap_4
XFILLER_61_127 VPWR VGND sg13g2_fill_2
X_12753_ net1864 fp16_res_pipe.x2\[5\] net1957 _00915_ VPWR VGND sg13g2_mux2_1
X_11704_ _05607_ VPWR _05608_ VGND _04585_ net1727 sg13g2_o21ai_1
X_14423_ _00224_ VGND VPWR _00962_ fpmul.seg_reg0.q\[8\] clknet_leaf_79_clk sg13g2_dfrbpq_1
X_12684_ _06495_ VPWR _00936_ VGND _06481_ _06494_ sg13g2_o21ai_1
XFILLER_24_70 VPWR VGND sg13g2_decap_8
X_11635_ net1837 VPWR _05540_ VGND _05435_ _05444_ sg13g2_o21ai_1
X_14354_ _00155_ VGND VPWR _00896_ _00007_ clknet_leaf_84_clk sg13g2_dfrbpq_1
XFILLER_11_783 VPWR VGND sg13g2_decap_8
X_13305_ acc\[2\] net1677 _07017_ VPWR VGND sg13g2_nor2_1
X_14285_ _00086_ VGND VPWR _07114_ fp16_sum_pipe.reg1en.d\[0\] clknet_leaf_53_clk
+ sg13g2_dfrbpq_2
X_10517_ _04559_ _04557_ _04558_ _04483_ net1737 VPWR VGND sg13g2_a22oi_1
X_13236_ _06961_ _02628_ _06960_ VPWR VGND sg13g2_nand2b_1
XFILLER_6_286 VPWR VGND sg13g2_decap_8
X_11497_ VPWR _05402_ fp16_sum_pipe.add_renorm0.mantisa\[5\] VGND sg13g2_inv_1
XFILLER_40_91 VPWR VGND sg13g2_decap_8
X_10448_ _04468_ _04496_ _04497_ VPWR VGND sg13g2_nor2_1
XFILLER_123_140 VPWR VGND sg13g2_decap_8
XFILLER_112_803 VPWR VGND sg13g2_decap_8
X_10379_ _04429_ _04423_ _04428_ VPWR VGND sg13g2_nand2_1
XFILLER_97_569 VPWR VGND sg13g2_decap_8
XFILLER_97_536 VPWR VGND sg13g2_fill_1
X_13098_ _06801_ _06790_ _06858_ VPWR VGND _06768_ sg13g2_nand3b_1
X_12118_ VGND VPWR _05956_ _05961_ _05964_ _05963_ sg13g2_a21oi_1
X_12049_ net1860 net1863 net1859 _05895_ VPWR VGND sg13g2_nand3_1
XFILLER_78_783 VPWR VGND sg13g2_fill_1
XFILLER_77_282 VPWR VGND sg13g2_fill_2
XFILLER_66_934 VPWR VGND sg13g2_fill_1
XFILLER_81_915 VPWR VGND sg13g2_decap_4
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_93_786 VPWR VGND sg13g2_decap_8
X_07590_ _01900_ _01903_ _01904_ VPWR VGND sg13g2_nor2_1
XFILLER_92_285 VPWR VGND sg13g2_fill_1
XFILLER_80_414 VPWR VGND sg13g2_fill_2
XFILLER_65_477 VPWR VGND sg13g2_fill_1
XFILLER_52_116 VPWR VGND sg13g2_decap_8
XFILLER_34_820 VPWR VGND sg13g2_fill_2
XFILLER_18_371 VPWR VGND sg13g2_decap_4
XFILLER_19_894 VPWR VGND sg13g2_decap_8
XFILLER_80_436 VPWR VGND sg13g2_fill_2
X_09260_ VPWR _03414_ fp16_res_pipe.op_sign_logic0.mantisa_b\[1\] VGND sg13g2_inv_1
XFILLER_61_694 VPWR VGND sg13g2_decap_4
XFILLER_60_182 VPWR VGND sg13g2_decap_8
X_08211_ _02467_ fp16_sum_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_inv_2
XFILLER_21_514 VPWR VGND sg13g2_decap_8
X_09191_ _03350_ VPWR _01283_ VGND net1906 _03349_ sg13g2_o21ai_1
XFILLER_21_569 VPWR VGND sg13g2_fill_2
X_08142_ _02403_ _02402_ _02352_ VPWR VGND sg13g2_nand2_1
XFILLER_107_619 VPWR VGND sg13g2_fill_2
XFILLER_107_608 VPWR VGND sg13g2_decap_8
XFILLER_106_107 VPWR VGND sg13g2_fill_2
Xplace1910 fp16_res_pipe.reg1en.d\[0\] net1910 VPWR VGND sg13g2_buf_2
XFILLER_20_28 VPWR VGND sg13g2_decap_8
Xplace1921 net1920 net1921 VPWR VGND sg13g2_buf_2
Xplace1943 net1941 net1943 VPWR VGND sg13g2_buf_2
Xplace1954 fpmul.reg1en.d\[0\] net1954 VPWR VGND sg13g2_buf_2
Xplace1932 net1930 net1932 VPWR VGND sg13g2_buf_1
XFILLER_114_140 VPWR VGND sg13g2_decap_8
XFILLER_0_407 VPWR VGND sg13g2_decap_8
X_08975_ VPWR _03161_ _03160_ VGND sg13g2_inv_1
XFILLER_103_869 VPWR VGND sg13g2_fill_2
XFILLER_69_772 VPWR VGND sg13g2_fill_1
XFILLER_69_761 VPWR VGND sg13g2_fill_1
XFILLER_29_603 VPWR VGND sg13g2_fill_1
X_07926_ _02198_ _02200_ _02201_ VPWR VGND sg13g2_nor2_1
XFILLER_111_880 VPWR VGND sg13g2_decap_8
XFILLER_68_282 VPWR VGND sg13g2_fill_2
XFILLER_68_271 VPWR VGND sg13g2_decap_8
XFILLER_57_945 VPWR VGND sg13g2_decap_8
XFILLER_56_422 VPWR VGND sg13g2_fill_1
X_07857_ _02151_ _02018_ net1795 VPWR VGND sg13g2_nand2_1
XFILLER_56_455 VPWR VGND sg13g2_decap_4
XFILLER_29_658 VPWR VGND sg13g2_decap_8
X_07788_ VPWR _02087_ acc_sub.exp_mant_logic0.b\[2\] VGND sg13g2_inv_1
XFILLER_83_285 VPWR VGND sg13g2_decap_8
XFILLER_45_14 VPWR VGND sg13g2_decap_8
XFILLER_43_105 VPWR VGND sg13g2_decap_8
X_09527_ _03644_ _03642_ _03643_ VPWR VGND sg13g2_nand2_1
XFILLER_72_959 VPWR VGND sg13g2_decap_4
XFILLER_43_149 VPWR VGND sg13g2_fill_1
XFILLER_24_330 VPWR VGND sg13g2_decap_8
XFILLER_25_831 VPWR VGND sg13g2_decap_4
XFILLER_101_42 VPWR VGND sg13g2_decap_8
XFILLER_101_20 VPWR VGND sg13g2_decap_8
XFILLER_71_469 VPWR VGND sg13g2_decap_4
XFILLER_40_812 VPWR VGND sg13g2_decap_8
XFILLER_24_352 VPWR VGND sg13g2_decap_8
XFILLER_61_13 VPWR VGND sg13g2_fill_1
XFILLER_52_694 VPWR VGND sg13g2_decap_8
X_09458_ _03590_ acc_sub.x2\[14\] net1915 VPWR VGND sg13g2_nand2_1
X_08409_ _02644_ fpdiv.divider0.counter\[3\] VPWR VGND sg13g2_inv_2
XFILLER_61_57 VPWR VGND sg13g2_fill_1
X_09389_ _03535_ _03492_ net1675 _03536_ VPWR VGND sg13g2_mux2_1
X_11420_ VGND VPWR _03327_ net1942 _01060_ _05356_ sg13g2_a21oi_1
XFILLER_125_405 VPWR VGND sg13g2_fill_2
X_11351_ VGND VPWR net1811 _05192_ _05304_ _05303_ sg13g2_a21oi_1
XFILLER_126_939 VPWR VGND sg13g2_decap_8
X_10302_ _04369_ net1911 fp16_res_pipe.x2\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_4_702 VPWR VGND sg13g2_decap_4
X_14070_ VPWR _00621_ net95 VGND sg13g2_inv_1
X_11282_ _05243_ acc_sum.exp_mant_logic0.a\[3\] _05192_ acc_sum.exp_mant_logic0.a\[2\]
+ net1653 VPWR VGND sg13g2_a22oi_1
XFILLER_3_223 VPWR VGND sg13g2_fill_1
XFILLER_79_525 VPWR VGND sg13g2_decap_8
XFILLER_79_514 VPWR VGND sg13g2_decap_8
X_10233_ _04304_ _04305_ _04297_ _04306_ VPWR VGND sg13g2_nand3_1
XFILLER_86_21 VPWR VGND sg13g2_fill_1
XFILLER_3_289 VPWR VGND sg13g2_fill_2
X_10164_ _04243_ VPWR _04244_ VGND _03607_ _04222_ sg13g2_o21ai_1
XFILLER_120_154 VPWR VGND sg13g2_decap_8
XFILLER_94_506 VPWR VGND sg13g2_decap_8
XFILLER_0_996 VPWR VGND sg13g2_decap_8
X_10095_ _04180_ _04179_ net1637 VPWR VGND sg13g2_nand2_1
XFILLER_19_113 VPWR VGND sg13g2_decap_8
XFILLER_75_764 VPWR VGND sg13g2_decap_8
XFILLER_74_241 VPWR VGND sg13g2_fill_2
XFILLER_74_230 VPWR VGND sg13g2_decap_4
X_13923_ VPWR _00474_ net11 VGND sg13g2_inv_1
XFILLER_19_70 VPWR VGND sg13g2_decap_4
XFILLER_74_252 VPWR VGND sg13g2_fill_2
XFILLER_63_948 VPWR VGND sg13g2_decap_8
XFILLER_63_915 VPWR VGND sg13g2_decap_8
X_13854_ VPWR _00405_ net29 VGND sg13g2_inv_1
XFILLER_35_639 VPWR VGND sg13g2_decap_8
XFILLER_34_105 VPWR VGND sg13g2_decap_8
XFILLER_19_168 VPWR VGND sg13g2_fill_2
XFILLER_90_745 VPWR VGND sg13g2_fill_1
XFILLER_16_820 VPWR VGND sg13g2_decap_8
XFILLER_28_691 VPWR VGND sg13g2_decap_8
X_13785_ VPWR _00336_ net126 VGND sg13g2_inv_1
XFILLER_15_363 VPWR VGND sg13g2_decap_8
XFILLER_16_875 VPWR VGND sg13g2_decap_8
X_10997_ _04984_ VPWR _01111_ VGND net1929 _02466_ sg13g2_o21ai_1
X_12736_ _06538_ VPWR _00927_ VGND _06536_ _02648_ sg13g2_o21ai_1
XFILLER_42_182 VPWR VGND sg13g2_decap_8
XFILLER_35_91 VPWR VGND sg13g2_decap_8
XFILLER_15_374 VPWR VGND sg13g2_fill_2
XFILLER_31_834 VPWR VGND sg13g2_decap_8
X_12667_ _06482_ _06415_ _06467_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_867 VPWR VGND sg13g2_fill_1
X_14406_ _00207_ VGND VPWR _00945_ fpmul.reg_a_out\[3\] clknet_leaf_100_clk sg13g2_dfrbpq_2
X_11618_ _05522_ VPWR _05523_ VGND _05517_ _05521_ sg13g2_o21ai_1
XFILLER_117_928 VPWR VGND sg13g2_decap_8
X_14337_ _00138_ VGND VPWR _00879_ fpmul.reg_p_out\[1\] clknet_leaf_82_clk sg13g2_dfrbpq_1
X_12598_ _06413_ _06411_ _06414_ VPWR VGND sg13g2_xor2_1
X_11549_ _05454_ _05452_ _05453_ VPWR VGND sg13g2_nand2_1
XFILLER_116_449 VPWR VGND sg13g2_fill_1
X_14268_ _00069_ VGND VPWR _00819_ fp16_res_pipe.x2\[1\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_14199_ VPWR _00750_ net105 VGND sg13g2_inv_1
XFILLER_97_300 VPWR VGND sg13g2_decap_8
X_13219_ _06946_ VPWR _06947_ VGND sipo.bit_counter\[2\] _06945_ sg13g2_o21ai_1
XFILLER_97_333 VPWR VGND sg13g2_decap_4
XFILLER_112_677 VPWR VGND sg13g2_fill_2
XFILLER_111_143 VPWR VGND sg13g2_fill_1
X_08760_ _02953_ acc_sum.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_inv_2
X_07711_ _01927_ net1660 _02018_ VPWR VGND sg13g2_nor2_2
X_08691_ net1817 acc_sum.add_renorm0.mantisa\[3\] _02906_ VPWR VGND sg13g2_nor2_1
XFILLER_18_0 VPWR VGND sg13g2_decap_8
X_07642_ _01953_ _01954_ _01952_ _01955_ VPWR VGND sg13g2_nand3_1
XFILLER_81_723 VPWR VGND sg13g2_decap_8
XFILLER_54_948 VPWR VGND sg13g2_decap_8
XFILLER_54_926 VPWR VGND sg13g2_fill_1
XFILLER_54_915 VPWR VGND sg13g2_decap_8
XFILLER_38_488 VPWR VGND sg13g2_decap_4
XFILLER_26_628 VPWR VGND sg13g2_fill_1
XFILLER_25_127 VPWR VGND sg13g2_fill_2
X_07573_ _01885_ _01886_ _01887_ VPWR VGND sg13g2_nor2b_1
X_09312_ _03465_ _03463_ _03464_ VPWR VGND sg13g2_nand2_1
XFILLER_15_28 VPWR VGND sg13g2_decap_8
XFILLER_40_119 VPWR VGND sg13g2_decap_8
XFILLER_34_694 VPWR VGND sg13g2_fill_2
XFILLER_22_812 VPWR VGND sg13g2_decap_8
X_09243_ _03397_ _03396_ VPWR VGND sg13g2_inv_2
XFILLER_21_355 VPWR VGND sg13g2_decap_8
XFILLER_119_210 VPWR VGND sg13g2_decap_8
X_09174_ _03339_ acc_sum.exp_mant_logic0.b\[9\] VPWR VGND sg13g2_inv_2
X_08125_ _02267_ _02349_ _02387_ VPWR VGND sg13g2_nor2_1
XFILLER_31_49 VPWR VGND sg13g2_decap_8
X_08056_ _02322_ _02307_ _02321_ VPWR VGND sg13g2_nand2_2
XFILLER_116_961 VPWR VGND sg13g2_decap_8
XFILLER_89_801 VPWR VGND sg13g2_decap_8
Xplace1740 _02726_ net1740 VPWR VGND sg13g2_buf_2
Xplace1762 net1761 net1762 VPWR VGND sg13g2_buf_2
Xplace1751 _06903_ net1751 VPWR VGND sg13g2_buf_2
Xplace1784 net1783 net1784 VPWR VGND sg13g2_buf_2
XFILLER_115_493 VPWR VGND sg13g2_fill_1
Xplace1773 _02965_ net1773 VPWR VGND sg13g2_buf_2
XFILLER_103_622 VPWR VGND sg13g2_decap_4
Xplace1795 acc_sub.exp_mant_logic0.b\[5\] net1795 VPWR VGND sg13g2_buf_2
X_08958_ _03144_ _01709_ _03143_ VPWR VGND sg13g2_xnor2_1
XFILLER_102_165 VPWR VGND sg13g2_decap_8
XFILLER_57_731 VPWR VGND sg13g2_fill_2
XFILLER_29_422 VPWR VGND sg13g2_fill_1
X_08889_ _03076_ _03062_ _03068_ VPWR VGND sg13g2_xnor2_1
XFILLER_91_509 VPWR VGND sg13g2_decap_8
XFILLER_56_230 VPWR VGND sg13g2_fill_1
XFILLER_45_904 VPWR VGND sg13g2_decap_4
X_07909_ _02184_ fp16_sum_pipe.exp_mant_logic0.a\[14\] fp16_sum_pipe.exp_mant_logic0.b\[14\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_84_583 VPWR VGND sg13g2_fill_2
XFILLER_57_797 VPWR VGND sg13g2_decap_4
XFILLER_56_274 VPWR VGND sg13g2_decap_8
XFILLER_56_252 VPWR VGND sg13g2_decap_8
XFILLER_44_414 VPWR VGND sg13g2_decap_8
X_10920_ _01132_ _04927_ _04928_ VPWR VGND sg13g2_nand2_1
XFILLER_17_617 VPWR VGND sg13g2_fill_1
XFILLER_29_488 VPWR VGND sg13g2_decap_8
XFILLER_56_296 VPWR VGND sg13g2_decap_8
XFILLER_56_285 VPWR VGND sg13g2_fill_2
XFILLER_45_948 VPWR VGND sg13g2_decap_8
XFILLER_16_138 VPWR VGND sg13g2_fill_2
XFILLER_112_63 VPWR VGND sg13g2_decap_8
XFILLER_72_778 VPWR VGND sg13g2_fill_1
XFILLER_72_767 VPWR VGND sg13g2_fill_1
XFILLER_72_34 VPWR VGND sg13g2_decap_8
XFILLER_60_929 VPWR VGND sg13g2_decap_8
X_10851_ net1824 fp16_res_pipe.add_renorm0.exp\[0\] _04863_ VPWR VGND sg13g2_nor2_1
XFILLER_53_981 VPWR VGND sg13g2_decap_8
X_13570_ VPWR _00121_ net27 VGND sg13g2_inv_1
XFILLER_25_683 VPWR VGND sg13g2_decap_8
X_10782_ VPWR _04794_ _04793_ VGND sg13g2_inv_1
X_12521_ _06346_ acc_sub.x2\[6\] VPWR VGND sg13g2_inv_2
XFILLER_13_856 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_fill_1
X_12452_ _00968_ _06295_ _06296_ VPWR VGND sg13g2_nand2_1
XFILLER_40_697 VPWR VGND sg13g2_fill_1
XFILLER_40_686 VPWR VGND sg13g2_decap_8
XFILLER_8_326 VPWR VGND sg13g2_fill_2
XFILLER_122_0 VPWR VGND sg13g2_decap_8
X_11403_ _05346_ VPWR _01067_ VGND _05345_ net1706 sg13g2_o21ai_1
XFILLER_8_348 VPWR VGND sg13g2_decap_8
XFILLER_126_736 VPWR VGND sg13g2_decap_8
X_12383_ _05891_ _06015_ _06225_ _06229_ VPWR VGND sg13g2_nor3_1
XFILLER_125_224 VPWR VGND sg13g2_decap_8
XFILLER_114_909 VPWR VGND sg13g2_decap_8
X_14122_ VPWR _00673_ net105 VGND sg13g2_inv_1
XFILLER_107_950 VPWR VGND sg13g2_decap_8
X_11334_ _03347_ _05148_ _05288_ VPWR VGND sg13g2_nor2_1
XFILLER_4_532 VPWR VGND sg13g2_decap_8
XFILLER_21_82 VPWR VGND sg13g2_fill_2
XFILLER_113_408 VPWR VGND sg13g2_fill_1
X_14053_ VPWR _00604_ net81 VGND sg13g2_inv_1
X_11265_ _05228_ _05073_ _05227_ net1808 _05211_ VPWR VGND sg13g2_a22oi_1
XFILLER_122_931 VPWR VGND sg13g2_decap_8
X_13004_ _06772_ fpmul.seg_reg0.q\[15\] fpmul.seg_reg0.q\[12\] VPWR VGND sg13g2_nand2_1
X_10216_ VGND VPWR fp16_res_pipe.exp_mant_logic0.b\[4\] net1644 _04290_ _04289_ sg13g2_a21oi_1
XFILLER_79_366 VPWR VGND sg13g2_decap_8
X_11196_ _05164_ _05162_ _05163_ VPWR VGND sg13g2_nand2_1
XFILLER_79_388 VPWR VGND sg13g2_decap_8
XFILLER_0_771 VPWR VGND sg13g2_decap_8
X_14955_ _00756_ VGND VPWR _01475_ acc_sub.add_renorm0.exp\[7\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_48_764 VPWR VGND sg13g2_fill_2
XFILLER_48_731 VPWR VGND sg13g2_fill_2
XFILLER_0_793 VPWR VGND sg13g2_decap_8
XFILLER_11_7 VPWR VGND sg13g2_decap_8
X_10078_ _04164_ net1827 net1643 net1688 fp16_res_pipe.exp_mant_logic0.a\[4\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_48_797 VPWR VGND sg13g2_fill_1
X_13906_ VPWR _00457_ net12 VGND sg13g2_inv_1
XFILLER_90_520 VPWR VGND sg13g2_decap_8
X_14886_ _00687_ VGND VPWR _01406_ acc_sub.exp_mant_logic0.b\[12\] clknet_leaf_55_clk
+ sg13g2_dfrbpq_2
XFILLER_63_745 VPWR VGND sg13g2_fill_2
XFILLER_47_296 VPWR VGND sg13g2_fill_1
XFILLER_36_948 VPWR VGND sg13g2_decap_8
XFILLER_51_907 VPWR VGND sg13g2_fill_2
X_13837_ VPWR _00388_ net14 VGND sg13g2_inv_1
X_13768_ VPWR _00319_ net109 VGND sg13g2_inv_1
XFILLER_22_108 VPWR VGND sg13g2_fill_1
X_12719_ _06478_ _06524_ _06523_ _06525_ VPWR VGND sg13g2_nand3_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
XFILLER_31_631 VPWR VGND sg13g2_decap_8
XFILLER_31_642 VPWR VGND sg13g2_fill_2
XFILLER_31_653 VPWR VGND sg13g2_fill_2
X_13699_ VPWR _00250_ net54 VGND sg13g2_inv_1
XFILLER_30_152 VPWR VGND sg13g2_fill_1
XFILLER_117_725 VPWR VGND sg13g2_decap_8
XFILLER_8_860 VPWR VGND sg13g2_decap_8
XFILLER_105_909 VPWR VGND sg13g2_decap_8
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_116_257 VPWR VGND sg13g2_decap_8
X_09930_ VPWR _04027_ _04026_ VGND sg13g2_inv_1
XFILLER_113_942 VPWR VGND sg13g2_decap_8
XFILLER_98_631 VPWR VGND sg13g2_decap_8
XFILLER_98_620 VPWR VGND sg13g2_fill_2
XFILLER_112_430 VPWR VGND sg13g2_decap_8
X_09861_ _03970_ _03968_ _03969_ _03967_ net1769 VPWR VGND sg13g2_a22oi_1
XFILLER_98_653 VPWR VGND sg13g2_fill_2
X_08812_ _02973_ _02991_ _02998_ _02999_ VPWR VGND sg13g2_nor3_2
X_09792_ VPWR _03906_ _03834_ VGND sg13g2_inv_1
XFILLER_100_636 VPWR VGND sg13g2_decap_8
XFILLER_86_848 VPWR VGND sg13g2_fill_2
XFILLER_100_669 VPWR VGND sg13g2_decap_8
XFILLER_100_647 VPWR VGND sg13g2_fill_2
X_08743_ _02942_ acc\[11\] net1901 VPWR VGND sg13g2_nand2_1
XFILLER_38_230 VPWR VGND sg13g2_decap_8
XFILLER_39_775 VPWR VGND sg13g2_decap_8
XFILLER_38_263 VPWR VGND sg13g2_fill_2
XFILLER_27_904 VPWR VGND sg13g2_decap_8
XFILLER_93_380 VPWR VGND sg13g2_fill_2
X_08674_ _02724_ VPWR _02891_ VGND _02850_ net1668 sg13g2_o21ai_1
XFILLER_66_583 VPWR VGND sg13g2_fill_1
XFILLER_53_211 VPWR VGND sg13g2_decap_8
X_07625_ VPWR _01939_ _01938_ VGND sg13g2_inv_1
XFILLER_81_564 VPWR VGND sg13g2_fill_1
XFILLER_26_49 VPWR VGND sg13g2_decap_8
XFILLER_26_469 VPWR VGND sg13g2_fill_1
X_07556_ _01870_ VPWR _01431_ VGND acc_sub.reg1en.q\[0\] _01499_ sg13g2_o21ai_1
XFILLER_35_981 VPWR VGND sg13g2_decap_8
X_07487_ _01807_ _01809_ _01810_ VPWR VGND sg13g2_nor2_2
X_09226_ VPWR _03380_ fp16_res_pipe.op_sign_logic0.mantisa_b\[7\] VGND sg13g2_inv_1
XFILLER_108_703 VPWR VGND sg13g2_decap_8
X_09157_ net1896 acc_sum.exp_mant_logic0.b\[15\] _03328_ VPWR VGND sg13g2_nor2_1
XFILLER_5_329 VPWR VGND sg13g2_decap_8
X_09088_ _03271_ VPWR _01307_ VGND net1801 _03259_ sg13g2_o21ai_1
X_08108_ _02371_ net1658 _02273_ VPWR VGND sg13g2_nand2_1
XFILLER_107_279 VPWR VGND sg13g2_decap_4
X_08039_ _02305_ _02294_ _02304_ VPWR VGND sg13g2_nand2_2
XFILLER_122_238 VPWR VGND sg13g2_decap_8
XFILLER_1_513 VPWR VGND sg13g2_decap_8
XFILLER_27_1002 VPWR VGND sg13g2_decap_8
XFILLER_104_964 VPWR VGND sg13g2_decap_8
X_11050_ _01102_ _04996_ _05028_ net1760 _04992_ VPWR VGND sg13g2_a22oi_1
XFILLER_27_1013 VPWR VGND sg13g2_fill_1
X_10001_ VGND VPWR _04078_ _04051_ _04089_ _04088_ sg13g2_a21oi_1
X_14740_ _00541_ VGND VPWR _01268_ fp16_res_pipe.add_renorm0.mantisa\[3\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_2
XFILLER_123_84 VPWR VGND sg13g2_decap_8
XFILLER_83_11 VPWR VGND sg13g2_fill_1
X_11952_ _05812_ net1883 fpmul.reg_b_out\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_17_425 VPWR VGND sg13g2_decap_8
XFILLER_18_948 VPWR VGND sg13g2_decap_8
XFILLER_29_296 VPWR VGND sg13g2_decap_4
X_11883_ _05771_ VPWR _01012_ VGND _02644_ _05767_ sg13g2_o21ai_1
XFILLER_60_715 VPWR VGND sg13g2_decap_4
XFILLER_44_244 VPWR VGND sg13g2_fill_2
XFILLER_33_918 VPWR VGND sg13g2_decap_8
X_14671_ _00472_ VGND VPWR _01199_ fp16_res_pipe.op_sign_logic0.mantisa_b\[8\] clknet_leaf_140_clk
+ sg13g2_dfrbpq_1
X_10903_ _04913_ _04912_ net1772 VPWR VGND sg13g2_nand2_1
X_13622_ VPWR _00173_ net65 VGND sg13g2_inv_1
X_10834_ _04836_ _04845_ _04846_ VPWR VGND sg13g2_nor2_1
X_13553_ VPWR _00104_ net87 VGND sg13g2_inv_1
XFILLER_60_759 VPWR VGND sg13g2_decap_8
XFILLER_16_93 VPWR VGND sg13g2_decap_8
X_12504_ fpmul.reg_a_out\[13\] net1951 _06336_ VPWR VGND sg13g2_nor2_1
XFILLER_40_461 VPWR VGND sg13g2_decap_8
XFILLER_8_112 VPWR VGND sg13g2_decap_8
XFILLER_9_613 VPWR VGND sg13g2_decap_8
X_10765_ fp16_res_pipe.add_renorm0.exp\[1\] fp16_res_pipe.add_renorm0.exp\[0\] fp16_res_pipe.add_renorm0.exp\[2\]
+ _04777_ VPWR VGND sg13g2_nand3_1
X_13484_ VPWR _00035_ net22 VGND sg13g2_inv_1
X_10696_ _04709_ net1826 fp16_res_pipe.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_13_697 VPWR VGND sg13g2_decap_8
X_12435_ _06275_ _06260_ _06261_ _06281_ VPWR VGND sg13g2_nor3_1
XFILLER_32_70 VPWR VGND sg13g2_decap_8
XFILLER_126_544 VPWR VGND sg13g2_fill_1
XFILLER_126_533 VPWR VGND sg13g2_decap_8
XFILLER_126_522 VPWR VGND sg13g2_decap_8
X_12366_ _06211_ _06204_ _06212_ VPWR VGND sg13g2_xor2_1
XFILLER_8_189 VPWR VGND sg13g2_decap_8
XFILLER_114_728 VPWR VGND sg13g2_fill_2
X_11317_ _05273_ net1697 acc_sum.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_59_7 VPWR VGND sg13g2_decap_4
XFILLER_4_351 VPWR VGND sg13g2_decap_8
X_14105_ VPWR _00656_ net42 VGND sg13g2_inv_1
XFILLER_113_216 VPWR VGND sg13g2_decap_8
X_12297_ VGND VPWR _06126_ _06132_ _06143_ _06142_ sg13g2_a21oi_1
XFILLER_5_885 VPWR VGND sg13g2_decap_8
X_14036_ VPWR _00587_ net99 VGND sg13g2_inv_1
XFILLER_80_1004 VPWR VGND sg13g2_decap_8
XFILLER_110_934 VPWR VGND sg13g2_decap_8
XFILLER_79_163 VPWR VGND sg13g2_decap_4
X_11179_ _05148_ _05146_ VPWR VGND sg13g2_inv_2
XFILLER_94_122 VPWR VGND sg13g2_decap_8
XFILLER_95_678 VPWR VGND sg13g2_decap_8
XFILLER_82_317 VPWR VGND sg13g2_decap_8
X_14938_ _00739_ VGND VPWR _01458_ acc_sub.exp_mant_logic0.a\[6\] clknet_leaf_56_clk
+ sg13g2_dfrbpq_2
XFILLER_82_328 VPWR VGND sg13g2_fill_1
XFILLER_36_778 VPWR VGND sg13g2_decap_8
X_14869_ _00670_ VGND VPWR _01393_ fp16_sum_pipe.op_sign_logic0.s_a clknet_leaf_112_clk
+ sg13g2_dfrbpq_1
XFILLER_24_918 VPWR VGND sg13g2_decap_8
X_07410_ _01748_ VPWR _01455_ VGND net1891 _01747_ sg13g2_o21ai_1
X_08390_ instr\[1\] _02612_ _02627_ VPWR VGND sg13g2_nor2_1
XFILLER_63_586 VPWR VGND sg13g2_fill_2
X_07341_ _01702_ net1665 _01586_ VPWR VGND sg13g2_nand2_1
XFILLER_85_0 VPWR VGND sg13g2_decap_8
X_07272_ _01507_ _01577_ _01504_ _01641_ VPWR VGND sg13g2_a21o_1
XFILLER_31_483 VPWR VGND sg13g2_decap_8
X_09011_ _03183_ _03196_ _03197_ VPWR VGND sg13g2_nor2_1
XFILLER_117_511 VPWR VGND sg13g2_fill_2
XFILLER_117_577 VPWR VGND sg13g2_fill_1
XFILLER_99_951 VPWR VGND sg13g2_decap_8
X_09913_ fp16_res_pipe.exp_mant_logic0.b\[8\] fp16_res_pipe.exp_mant_logic0.a\[8\]
+ _04010_ VPWR VGND sg13g2_xor2_1
XFILLER_101_934 VPWR VGND sg13g2_decap_8
X_09844_ _03952_ _03954_ _03783_ _03955_ VPWR VGND sg13g2_nand3_1
XFILLER_86_645 VPWR VGND sg13g2_fill_1
X_09775_ _03890_ _03861_ _03867_ VPWR VGND sg13g2_nand2_1
XFILLER_85_177 VPWR VGND sg13g2_decap_8
XFILLER_67_870 VPWR VGND sg13g2_fill_2
XFILLER_96_1011 VPWR VGND sg13g2_fill_2
X_08726_ _02931_ net1815 acc_sum.seg_reg0.q\[23\] VPWR VGND sg13g2_nand2_1
XFILLER_26_211 VPWR VGND sg13g2_decap_8
X_08657_ VPWR _02876_ _02852_ VGND sg13g2_inv_1
X_07608_ _01910_ _01921_ _01922_ VPWR VGND sg13g2_nor2_1
XFILLER_53_14 VPWR VGND sg13g2_decap_8
XFILLER_27_789 VPWR VGND sg13g2_decap_8
X_08588_ _02811_ acc_sum.op_sign_logic0.mantisa_a\[8\] acc_sum.op_sign_logic0.mantisa_b\[8\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_23_940 VPWR VGND sg13g2_decap_8
X_07539_ _01857_ _01844_ acc_sub.exp_mant_logic0.b\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_41_258 VPWR VGND sg13g2_decap_8
XFILLER_50_792 VPWR VGND sg13g2_decap_8
X_10550_ _04585_ fp16_sum_pipe.add_renorm0.exp\[5\] VPWR VGND sg13g2_inv_2
XFILLER_22_483 VPWR VGND sg13g2_decap_8
XFILLER_127_308 VPWR VGND sg13g2_decap_8
X_09209_ _03364_ fp16_res_pipe.op_sign_logic0.add_sub _03363_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_667 VPWR VGND sg13g2_fill_2
X_10481_ _04528_ _04397_ _04527_ VPWR VGND sg13g2_xnor2_1
XFILLER_108_522 VPWR VGND sg13g2_decap_8
X_12220_ _06066_ _06064_ _06065_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_126 VPWR VGND sg13g2_decap_8
XFILLER_108_555 VPWR VGND sg13g2_decap_8
XFILLER_2_800 VPWR VGND sg13g2_decap_8
XFILLER_123_525 VPWR VGND sg13g2_fill_2
XFILLER_123_514 VPWR VGND sg13g2_decap_8
XFILLER_118_84 VPWR VGND sg13g2_decap_8
XFILLER_78_11 VPWR VGND sg13g2_fill_2
X_12151_ VPWR _05997_ _05995_ VGND sg13g2_inv_1
X_11102_ _05072_ _05073_ VPWR VGND sg13g2_inv_4
X_12082_ _05928_ _05924_ _05927_ VPWR VGND sg13g2_nand2_1
XFILLER_103_260 VPWR VGND sg13g2_decap_4
XFILLER_76_100 VPWR VGND sg13g2_decap_8
X_11033_ acc_sum.exp_mant_logic0.b\[10\] _02943_ _05012_ VPWR VGND sg13g2_nor2_1
XFILLER_2_877 VPWR VGND sg13g2_decap_8
XFILLER_76_133 VPWR VGND sg13g2_fill_2
XFILLER_1_387 VPWR VGND sg13g2_decap_8
XFILLER_94_54 VPWR VGND sg13g2_decap_4
XFILLER_94_21 VPWR VGND sg13g2_decap_8
XFILLER_65_829 VPWR VGND sg13g2_decap_8
XFILLER_92_637 VPWR VGND sg13g2_fill_1
XFILLER_91_136 VPWR VGND sg13g2_decap_8
X_12984_ _06752_ _06751_ fpmul.seg_reg0.q\[18\] VPWR VGND sg13g2_nand2_1
XFILLER_45_520 VPWR VGND sg13g2_fill_2
XFILLER_18_745 VPWR VGND sg13g2_fill_1
XFILLER_94_98 VPWR VGND sg13g2_decap_8
X_11935_ _05800_ VPWR _00989_ VGND net1879 _05799_ sg13g2_o21ai_1
X_14723_ _00524_ VGND VPWR _01251_ fp16_res_pipe.exp_mant_logic0.a\[10\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
XFILLER_18_778 VPWR VGND sg13g2_decap_8
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_72_383 VPWR VGND sg13g2_fill_1
XFILLER_17_277 VPWR VGND sg13g2_fill_2
X_14654_ _00455_ VGND VPWR _01182_ fp16_res_pipe.exp_mant_logic0.b\[7\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_1
X_13605_ VPWR _00156_ net123 VGND sg13g2_inv_1
X_11866_ _05762_ net1756 add_result\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_14_951 VPWR VGND sg13g2_decap_8
X_11797_ net1837 _05698_ _05694_ _05699_ VPWR VGND sg13g2_nand3_1
X_14585_ _00386_ VGND VPWR _01117_ fp16_sum_pipe.exp_mant_logic0.b\[12\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_2
X_10817_ VPWR _04829_ _04828_ VGND sg13g2_inv_1
X_13536_ VPWR _00087_ net84 VGND sg13g2_inv_1
XFILLER_43_91 VPWR VGND sg13g2_decap_8
X_10748_ _04689_ _04690_ _04761_ VPWR VGND sg13g2_nor2_1
XFILLER_118_319 VPWR VGND sg13g2_decap_8
X_13467_ _02571_ _02564_ _00002_ VPWR VGND sg13g2_and2_1
XFILLER_9_465 VPWR VGND sg13g2_decap_8
XFILLER_127_820 VPWR VGND sg13g2_decap_8
X_12418_ _06263_ _06253_ _06264_ VPWR VGND sg13g2_xor2_1
X_10679_ _04647_ _04658_ _04692_ VPWR VGND sg13g2_nor2_1
X_13398_ VGND VPWR _06941_ _07055_ _00802_ _07075_ sg13g2_a21oi_1
XFILLER_127_897 VPWR VGND sg13g2_decap_8
XFILLER_126_374 VPWR VGND sg13g2_fill_1
X_12349_ _06195_ _06190_ _06194_ VPWR VGND sg13g2_xnor2_1
XFILLER_87_409 VPWR VGND sg13g2_decap_8
XFILLER_101_219 VPWR VGND sg13g2_fill_1
X_14019_ VPWR _00570_ net22 VGND sg13g2_inv_1
XFILLER_4_63 VPWR VGND sg13g2_decap_8
XFILLER_122_591 VPWR VGND sg13g2_decap_4
XFILLER_122_580 VPWR VGND sg13g2_fill_1
X_07890_ _02172_ net1892 acc_sub.x2\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_96_976 VPWR VGND sg13g2_decap_8
XFILLER_83_604 VPWR VGND sg13g2_fill_1
XFILLER_67_144 VPWR VGND sg13g2_fill_1
XFILLER_55_306 VPWR VGND sg13g2_decap_8
X_09560_ _03677_ _03659_ _03676_ VPWR VGND sg13g2_nand2_1
X_08511_ acc_sum.op_sign_logic0.mantisa_a\[7\] _02734_ _02735_ VPWR VGND sg13g2_nor2_1
XFILLER_70_309 VPWR VGND sg13g2_decap_4
X_09491_ _03612_ acc_sub.x2\[3\] net1918 VPWR VGND sg13g2_nand2_1
X_08442_ _02676_ _02674_ _02675_ VPWR VGND sg13g2_nand2_1
XFILLER_91_670 VPWR VGND sg13g2_decap_8
XFILLER_64_873 VPWR VGND sg13g2_decap_8
XFILLER_51_512 VPWR VGND sg13g2_decap_8
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_23_225 VPWR VGND sg13g2_fill_1
X_08373_ _02605_ _02615_ _02589_ _02616_ VPWR VGND sg13g2_nor3_1
XFILLER_23_28 VPWR VGND sg13g2_decap_8
X_07324_ _01686_ VPWR _01687_ VGND net1666 _01685_ sg13g2_o21ai_1
X_07255_ VPWR _01625_ _01624_ VGND sg13g2_inv_1
XFILLER_20_976 VPWR VGND sg13g2_decap_8
XFILLER_118_831 VPWR VGND sg13g2_decap_8
X_07186_ _01555_ _01557_ _01558_ VPWR VGND sg13g2_nor2_1
XFILLER_3_608 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_113_580 VPWR VGND sg13g2_fill_2
XFILLER_87_965 VPWR VGND sg13g2_decap_8
XFILLER_58_111 VPWR VGND sg13g2_decap_4
X_09827_ _03858_ _03880_ _03939_ VPWR VGND sg13g2_nor2_1
XFILLER_101_764 VPWR VGND sg13g2_decap_4
XFILLER_86_464 VPWR VGND sg13g2_fill_2
X_09758_ _03874_ _03873_ _03867_ VPWR VGND sg13g2_nand2_1
XFILLER_104_31 VPWR VGND sg13g2_decap_8
XFILLER_58_188 VPWR VGND sg13g2_decap_4
X_08709_ _02920_ acc_sum.add_renorm0.exp\[7\] VPWR VGND sg13g2_inv_2
XFILLER_64_35 VPWR VGND sg13g2_fill_1
X_09689_ acc_sum.add_renorm0.mantisa\[11\] acc_sum.add_renorm0.exp\[0\] _03805_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_73_169 VPWR VGND sg13g2_decap_8
XFILLER_55_873 VPWR VGND sg13g2_decap_8
X_11720_ _05608_ _05622_ _05624_ VPWR VGND sg13g2_nor2_1
XFILLER_42_545 VPWR VGND sg13g2_fill_2
XFILLER_120_63 VPWR VGND sg13g2_decap_8
XFILLER_70_887 VPWR VGND sg13g2_decap_4
XFILLER_42_578 VPWR VGND sg13g2_decap_8
Xfanout40 net41 net40 VPWR VGND sg13g2_buf_2
XFILLER_11_910 VPWR VGND sg13g2_decap_8
X_11651_ _05556_ _05477_ _05465_ _05428_ _05442_ VPWR VGND sg13g2_a22oi_1
XFILLER_30_718 VPWR VGND sg13g2_decap_4
Xfanout73 net74 net73 VPWR VGND sg13g2_buf_2
Xfanout62 net71 net62 VPWR VGND sg13g2_buf_2
Xfanout51 net56 net51 VPWR VGND sg13g2_buf_2
X_14370_ _00171_ VGND VPWR _00911_ fpmul.reg_b_out\[1\] clknet_leaf_106_clk sg13g2_dfrbpq_2
X_10602_ _04614_ VPWR _04615_ VGND fp16_res_pipe.add_renorm0.mantisa\[11\] _04613_
+ sg13g2_o21ai_1
XFILLER_10_420 VPWR VGND sg13g2_fill_1
X_11582_ _05469_ _05486_ _05487_ VPWR VGND sg13g2_nor2_1
XFILLER_127_105 VPWR VGND sg13g2_decap_8
Xfanout95 net96 net95 VPWR VGND sg13g2_buf_1
Xfanout84 net85 net84 VPWR VGND sg13g2_buf_2
XFILLER_6_402 VPWR VGND sg13g2_fill_1
X_10533_ net1849 fp16_sum_pipe.add_renorm0.mantisa\[2\] _04573_ VPWR VGND sg13g2_nor2_1
XFILLER_109_842 VPWR VGND sg13g2_decap_8
XFILLER_7_958 VPWR VGND sg13g2_decap_8
XFILLER_10_464 VPWR VGND sg13g2_fill_2
XFILLER_11_987 VPWR VGND sg13g2_decap_8
X_13252_ acc\[14\] _06975_ net1676 _00848_ VPWR VGND sg13g2_mux2_1
X_10464_ VPWR _04512_ _04511_ VGND sg13g2_inv_1
XFILLER_6_446 VPWR VGND sg13g2_decap_8
XFILLER_124_823 VPWR VGND sg13g2_decap_8
XFILLER_109_886 VPWR VGND sg13g2_decap_8
XFILLER_108_363 VPWR VGND sg13g2_decap_8
X_12203_ _06049_ _06046_ _06048_ VPWR VGND sg13g2_nand2_1
X_13183_ VPWR _06923_ sipo.shift_reg\[10\] VGND sg13g2_inv_1
X_10395_ _04445_ _04431_ _04444_ VPWR VGND sg13g2_nand2_1
X_12134_ VGND VPWR _05932_ _05936_ _05980_ _05979_ sg13g2_a21oi_1
XFILLER_96_228 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_104_591 VPWR VGND sg13g2_decap_8
X_12065_ VPWR _05911_ _05910_ VGND sg13g2_inv_1
XFILLER_49_133 VPWR VGND sg13g2_decap_8
XFILLER_77_497 VPWR VGND sg13g2_decap_8
XFILLER_64_125 VPWR VGND sg13g2_decap_8
XFILLER_93_968 VPWR VGND sg13g2_decap_8
Xclkbuf_5_24__f_clk clknet_4_12_0_clk clknet_5_24__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_65_659 VPWR VGND sg13g2_decap_4
XFILLER_64_158 VPWR VGND sg13g2_decap_8
XFILLER_38_91 VPWR VGND sg13g2_decap_8
X_12967_ _00006_ net1731 net1702 _06737_ VPWR VGND sg13g2_nand3_1
XFILLER_52_309 VPWR VGND sg13g2_decap_8
XFILLER_45_372 VPWR VGND sg13g2_decap_8
XFILLER_18_564 VPWR VGND sg13g2_decap_4
X_14706_ _00507_ VGND VPWR _01234_ acc_sum.y\[9\] clknet_leaf_48_clk sg13g2_dfrbpq_1
XFILLER_72_191 VPWR VGND sg13g2_fill_1
XFILLER_72_180 VPWR VGND sg13g2_decap_8
X_12898_ _06674_ net1910 fp16_res_pipe.y\[6\] VPWR VGND sg13g2_nand2_1
X_11918_ VPWR _05789_ fpmul.seg_reg0.q\[40\] VGND sg13g2_inv_1
X_14637_ _00438_ VGND VPWR _01169_ fp16_sum_pipe.add_renorm0.mantisa\[8\] clknet_leaf_109_clk
+ sg13g2_dfrbpq_1
XFILLER_21_718 VPWR VGND sg13g2_decap_8
X_11849_ _05747_ _05496_ _05617_ VPWR VGND sg13g2_nand2_1
XFILLER_33_578 VPWR VGND sg13g2_fill_1
X_14568_ _00369_ VGND VPWR _01104_ acc_sum.op_sign_logic0.s_a clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_20_239 VPWR VGND sg13g2_fill_1
XFILLER_118_105 VPWR VGND sg13g2_decap_8
Xclkload10 clknet_5_21__leaf_clk clkload10/Y VPWR VGND sg13g2_inv_4
X_14499_ _00300_ VGND VPWR _01035_ fpdiv.divider0.divisor\[10\] clknet_leaf_84_clk
+ sg13g2_dfrbpq_1
X_13519_ VPWR _00070_ net82 VGND sg13g2_inv_1
XFILLER_127_661 VPWR VGND sg13g2_decap_8
XFILLER_127_650 VPWR VGND sg13g2_decap_8
Xclkload32 clknet_leaf_10_clk clkload32/Y VPWR VGND sg13g2_inv_4
Xclkload21 VPWR clkload21/Y clknet_leaf_2_clk VGND sg13g2_inv_1
Xclkload43 clknet_leaf_135_clk clkload43/Y VPWR VGND sg13g2_inv_4
XFILLER_127_672 VPWR VGND sg13g2_decap_8
XFILLER_115_823 VPWR VGND sg13g2_decap_8
Xclkload87 clkload87/Y clknet_leaf_40_clk VPWR VGND sg13g2_inv_8
Xclkload76 clkload76/Y clknet_leaf_23_clk VPWR VGND sg13g2_inv_2
Xclkload65 clknet_leaf_101_clk clkload65/Y VPWR VGND sg13g2_inv_4
Xclkload54 clknet_leaf_93_clk clkload54/Y VPWR VGND sg13g2_inv_4
XFILLER_126_182 VPWR VGND sg13g2_decap_8
Xclkload98 clknet_leaf_79_clk clkload98/Y VPWR VGND sg13g2_inv_4
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_08991_ _03177_ _03167_ _03176_ VPWR VGND sg13g2_nand2_1
XFILLER_114_388 VPWR VGND sg13g2_decap_8
XFILLER_69_943 VPWR VGND sg13g2_decap_4
XFILLER_68_431 VPWR VGND sg13g2_decap_8
X_07942_ fp16_sum_pipe.exp_mant_logic0.a\[7\] _02216_ _02217_ VPWR VGND sg13g2_nor2_2
X_07873_ _02163_ VPWR _01407_ VGND net1889 _01784_ sg13g2_o21ai_1
XFILLER_84_924 VPWR VGND sg13g2_decap_8
X_09612_ _03726_ _03728_ _03729_ VPWR VGND sg13g2_nor2_1
XFILLER_18_28 VPWR VGND sg13g2_decap_8
X_09543_ VPWR _03660_ _03659_ VGND sg13g2_inv_1
XFILLER_93_1003 VPWR VGND sg13g2_decap_8
XFILLER_83_489 VPWR VGND sg13g2_fill_1
XFILLER_83_478 VPWR VGND sg13g2_decap_8
XFILLER_70_128 VPWR VGND sg13g2_fill_1
XFILLER_52_832 VPWR VGND sg13g2_decap_4
XFILLER_36_394 VPWR VGND sg13g2_fill_2
X_09474_ _03600_ VPWR _01250_ VGND net1920 _03599_ sg13g2_o21ai_1
X_08425_ _02659_ fpdiv.divider0.divisor_reg\[6\] fpdiv.divider0.remainder_reg\[6\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_54_1009 VPWR VGND sg13g2_decap_4
XFILLER_51_353 VPWR VGND sg13g2_decap_4
XFILLER_34_49 VPWR VGND sg13g2_decap_8
X_08356_ _02599_ _02598_ VPWR VGND sg13g2_inv_2
XFILLER_52_898 VPWR VGND sg13g2_decap_4
X_07307_ _01538_ _01671_ net1667 _01672_ VPWR VGND sg13g2_nor3_1
Xclkload4 VPWR clkload4/Y clknet_5_9__leaf_clk VGND sg13g2_inv_1
XFILLER_126_7 VPWR VGND sg13g2_decap_8
X_08287_ _02458_ _02427_ _02535_ VPWR VGND sg13g2_nor2_1
XFILLER_20_784 VPWR VGND sg13g2_decap_8
X_07238_ _01608_ VPWR _01609_ VGND _01523_ _01525_ sg13g2_o21ai_1
X_07169_ _01538_ _01540_ _01541_ VPWR VGND sg13g2_nor2_2
XFILLER_124_119 VPWR VGND sg13g2_decap_8
XFILLER_105_311 VPWR VGND sg13g2_decap_8
XFILLER_3_427 VPWR VGND sg13g2_decap_8
XFILLER_117_182 VPWR VGND sg13g2_decap_8
XFILLER_121_826 VPWR VGND sg13g2_decap_8
XFILLER_106_878 VPWR VGND sg13g2_fill_2
XFILLER_59_35 VPWR VGND sg13g2_decap_8
X_10180_ _03617_ _04233_ _04259_ VPWR VGND sg13g2_nor2_1
XFILLER_120_347 VPWR VGND sg13g2_decap_8
XFILLER_120_325 VPWR VGND sg13g2_fill_2
XFILLER_78_239 VPWR VGND sg13g2_fill_1
XFILLER_59_79 VPWR VGND sg13g2_decap_4
XFILLER_115_63 VPWR VGND sg13g2_decap_8
XFILLER_87_751 VPWR VGND sg13g2_decap_8
XFILLER_59_442 VPWR VGND sg13g2_decap_8
X_13870_ VPWR _00421_ net50 VGND sg13g2_inv_1
XFILLER_19_339 VPWR VGND sg13g2_decap_4
XFILLER_75_89 VPWR VGND sg13g2_fill_1
XFILLER_75_78 VPWR VGND sg13g2_decap_8
X_12821_ _06602_ _06603_ _06592_ _00907_ VPWR VGND sg13g2_nand3_1
XFILLER_74_456 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_fill_1
XFILLER_28_840 VPWR VGND sg13g2_decap_4
XFILLER_74_489 VPWR VGND sg13g2_decap_8
XFILLER_62_618 VPWR VGND sg13g2_decap_8
XFILLER_43_821 VPWR VGND sg13g2_fill_1
XFILLER_55_681 VPWR VGND sg13g2_decap_8
X_12752_ _06543_ VPWR _00916_ VGND net1956 _06031_ sg13g2_o21ai_1
XFILLER_43_832 VPWR VGND sg13g2_decap_8
X_12683_ _06495_ _06354_ div_result\[10\] VPWR VGND sg13g2_nand2_1
X_11703_ _05607_ net1727 _05606_ VPWR VGND sg13g2_nand2_1
X_14422_ _00223_ VGND VPWR _00961_ fpmul.seg_reg0.q\[7\] clknet_leaf_79_clk sg13g2_dfrbpq_1
XFILLER_70_684 VPWR VGND sg13g2_decap_8
X_11634_ _05534_ _05537_ _05533_ _05539_ VPWR VGND _05538_ sg13g2_nand4_1
XFILLER_11_751 VPWR VGND sg13g2_decap_8
X_14353_ _00154_ VGND VPWR _00895_ _00006_ clknet_leaf_82_clk sg13g2_dfrbpq_1
XFILLER_7_733 VPWR VGND sg13g2_fill_1
XFILLER_7_722 VPWR VGND sg13g2_decap_8
X_11565_ _05470_ fp16_sum_pipe.add_renorm0.mantisa\[4\] _05426_ VPWR VGND sg13g2_xnor2_1
X_13304_ VPWR VGND acc_sub.y\[2\] _07015_ _02578_ net1728 _07016_ acc_sum.y\[2\] sg13g2_a221oi_1
X_14284_ _00085_ VGND VPWR _07115_ fpdiv.reg1en.d\[0\] clknet_leaf_53_clk sg13g2_dfrbpq_2
X_10516_ VGND VPWR net1670 _04510_ _04558_ net1737 sg13g2_a21oi_1
X_11496_ VPWR _05401_ _05400_ VGND sg13g2_inv_1
XFILLER_124_620 VPWR VGND sg13g2_decap_8
XFILLER_115_119 VPWR VGND sg13g2_decap_8
XFILLER_109_694 VPWR VGND sg13g2_fill_1
XFILLER_108_160 VPWR VGND sg13g2_fill_2
X_13235_ _06960_ net1742 sipo.word_ready VPWR VGND sg13g2_nand2_1
XFILLER_40_70 VPWR VGND sg13g2_decap_8
X_10447_ _04496_ _04451_ _04495_ _04470_ _04386_ VPWR VGND sg13g2_a22oi_1
XFILLER_124_653 VPWR VGND sg13g2_decap_4
XFILLER_108_193 VPWR VGND sg13g2_decap_8
XFILLER_124_686 VPWR VGND sg13g2_fill_1
X_13166_ VPWR _06911_ sipo.shift_reg\[15\] VGND sg13g2_inv_1
XFILLER_41_7 VPWR VGND sg13g2_decap_8
X_10378_ _04425_ _04427_ _04428_ VPWR VGND sg13g2_nor2_2
XFILLER_123_196 VPWR VGND sg13g2_decap_8
XFILLER_112_859 VPWR VGND sg13g2_decap_8
XFILLER_111_314 VPWR VGND sg13g2_decap_8
XFILLER_97_548 VPWR VGND sg13g2_decap_8
X_13097_ _06768_ VPWR _06857_ VGND _06791_ _06856_ sg13g2_o21ai_1
X_12117_ VPWR _05963_ _05962_ VGND sg13g2_inv_1
XFILLER_3_994 VPWR VGND sg13g2_decap_8
XFILLER_2_493 VPWR VGND sg13g2_decap_8
XFILLER_78_751 VPWR VGND sg13g2_fill_1
X_12048_ VPWR _05894_ _05893_ VGND sg13g2_inv_1
XFILLER_93_732 VPWR VGND sg13g2_fill_1
XFILLER_93_743 VPWR VGND sg13g2_fill_2
XFILLER_66_957 VPWR VGND sg13g2_decap_4
XFILLER_65_445 VPWR VGND sg13g2_fill_2
XFILLER_65_434 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
X_13999_ VPWR _00550_ net30 VGND sg13g2_inv_1
XFILLER_18_350 VPWR VGND sg13g2_fill_2
XFILLER_25_309 VPWR VGND sg13g2_decap_8
XFILLER_74_990 VPWR VGND sg13g2_decap_4
XFILLER_60_172 VPWR VGND sg13g2_decap_8
XFILLER_34_898 VPWR VGND sg13g2_decap_8
X_08210_ _02466_ fp16_sum_pipe.exp_mant_logic0.b\[6\] VPWR VGND sg13g2_inv_2
X_09190_ _03350_ acc_sub.x2\[4\] net1906 VPWR VGND sg13g2_nand2_1
X_08141_ _02400_ _02401_ _02395_ _02402_ VPWR VGND sg13g2_nand3_1
Xclkload110 clkload110/Y clknet_leaf_72_clk VPWR VGND sg13g2_inv_2
X_08072_ _02305_ _02337_ _02338_ VPWR VGND sg13g2_nor2b_2
XFILLER_106_119 VPWR VGND sg13g2_fill_2
Xplace1900 net1897 net1900 VPWR VGND sg13g2_buf_2
Xplace1911 net1910 net1911 VPWR VGND sg13g2_buf_2
XFILLER_115_620 VPWR VGND sg13g2_fill_1
Xplace1944 fpdiv.reg1en.d\[0\] net1944 VPWR VGND sg13g2_buf_2
Xplace1922 fp16_sum_pipe.reg1en.d\[0\] net1922 VPWR VGND sg13g2_buf_1
Xplace1955 net1954 net1955 VPWR VGND sg13g2_buf_2
Xplace1933 net1930 net1933 VPWR VGND sg13g2_buf_2
XFILLER_115_686 VPWR VGND sg13g2_decap_8
X_08974_ _03160_ _01721_ _03159_ VPWR VGND sg13g2_xnor2_1
XFILLER_102_325 VPWR VGND sg13g2_decap_8
XFILLER_102_358 VPWR VGND sg13g2_decap_8
XFILLER_60_1013 VPWR VGND sg13g2_fill_1
XFILLER_60_1002 VPWR VGND sg13g2_decap_8
X_07925_ fp16_sum_pipe.exp_mant_logic0.a\[12\] _02199_ _02200_ VPWR VGND sg13g2_nor2_2
XFILLER_29_49 VPWR VGND sg13g2_decap_8
XFILLER_96_581 VPWR VGND sg13g2_fill_2
XFILLER_96_570 VPWR VGND sg13g2_decap_8
XFILLER_21_1008 VPWR VGND sg13g2_decap_4
X_07856_ _02150_ _02006_ acc_sub.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_84_765 VPWR VGND sg13g2_decap_8
XFILLER_84_743 VPWR VGND sg13g2_decap_8
XFILLER_57_968 VPWR VGND sg13g2_fill_1
XFILLER_28_147 VPWR VGND sg13g2_decap_8
X_07787_ _01416_ _02085_ _02086_ VPWR VGND sg13g2_nand2_1
XFILLER_72_927 VPWR VGND sg13g2_decap_4
XFILLER_28_158 VPWR VGND sg13g2_fill_2
X_09526_ _03643_ _03625_ _03619_ VPWR VGND sg13g2_nand2_1
XFILLER_71_448 VPWR VGND sg13g2_decap_8
XFILLER_52_651 VPWR VGND sg13g2_fill_2
X_09457_ VPWR _03589_ fp16_res_pipe.exp_mant_logic0.a\[14\] VGND sg13g2_inv_1
XFILLER_36_191 VPWR VGND sg13g2_decap_8
X_08408_ VPWR _02643_ fpdiv.divider0.state VGND sg13g2_inv_1
XFILLER_101_98 VPWR VGND sg13g2_decap_4
XFILLER_40_868 VPWR VGND sg13g2_decap_8
X_09388_ VGND VPWR _03420_ _03425_ _03535_ _03424_ sg13g2_a21oi_1
X_08339_ sipo.word\[14\] sipo.word\[13\] sipo.word\[15\] _02584_ VPWR VGND sipo.word\[12\]
+ sg13g2_nand4_1
XFILLER_126_918 VPWR VGND sg13g2_decap_8
X_11350_ _05303_ _05301_ _05302_ VPWR VGND sg13g2_nand2_1
XFILLER_4_725 VPWR VGND sg13g2_decap_8
X_10301_ _01191_ _04367_ _04368_ VPWR VGND sg13g2_nand2_1
X_13020_ _06784_ _06787_ _06781_ _06788_ VPWR VGND sg13g2_nand3_1
X_11281_ _05242_ net1809 _05227_ net1810 _05211_ VPWR VGND sg13g2_a22oi_1
XFILLER_4_747 VPWR VGND sg13g2_decap_8
XFILLER_4_769 VPWR VGND sg13g2_decap_8
XFILLER_3_257 VPWR VGND sg13g2_decap_8
X_10232_ _04305_ _04165_ net1830 VPWR VGND sg13g2_nand2_1
XFILLER_105_163 VPWR VGND sg13g2_fill_1
XFILLER_79_548 VPWR VGND sg13g2_decap_8
XFILLER_10_84 VPWR VGND sg13g2_decap_8
X_10163_ _04243_ _04224_ net1827 VPWR VGND sg13g2_nand2_1
XFILLER_126_84 VPWR VGND sg13g2_decap_8
XFILLER_120_133 VPWR VGND sg13g2_decap_8
XFILLER_86_33 VPWR VGND sg13g2_decap_8
XFILLER_48_902 VPWR VGND sg13g2_fill_2
XFILLER_0_975 VPWR VGND sg13g2_decap_8
XFILLER_86_66 VPWR VGND sg13g2_fill_1
XFILLER_75_710 VPWR VGND sg13g2_decap_8
X_10094_ _04173_ _04174_ _04172_ _04179_ VPWR VGND _04178_ sg13g2_nand4_1
XFILLER_75_754 VPWR VGND sg13g2_fill_2
XFILLER_59_283 VPWR VGND sg13g2_decap_8
XFILLER_48_979 VPWR VGND sg13g2_fill_1
XFILLER_48_957 VPWR VGND sg13g2_decap_8
X_13922_ VPWR _00473_ net5 VGND sg13g2_inv_1
XFILLER_90_702 VPWR VGND sg13g2_decap_8
XFILLER_74_264 VPWR VGND sg13g2_decap_8
XFILLER_62_404 VPWR VGND sg13g2_decap_8
X_13853_ VPWR _00404_ net30 VGND sg13g2_inv_1
XFILLER_16_810 VPWR VGND sg13g2_fill_1
XFILLER_90_757 VPWR VGND sg13g2_fill_2
XFILLER_74_297 VPWR VGND sg13g2_decap_8
X_12804_ _06587_ VPWR _06588_ VGND net1958 _06585_ sg13g2_o21ai_1
XFILLER_62_448 VPWR VGND sg13g2_fill_2
XFILLER_62_437 VPWR VGND sg13g2_decap_8
XFILLER_56_990 VPWR VGND sg13g2_decap_8
X_13784_ VPWR _00335_ net126 VGND sg13g2_inv_1
XFILLER_35_70 VPWR VGND sg13g2_decap_8
XFILLER_16_854 VPWR VGND sg13g2_decap_8
X_10996_ _04984_ fp16_res_pipe.x2\[6\] net1928 VPWR VGND sg13g2_nand2_1
X_12735_ _06513_ VPWR _06538_ VGND net1734 _06537_ sg13g2_o21ai_1
XFILLER_30_312 VPWR VGND sg13g2_fill_1
XFILLER_31_813 VPWR VGND sg13g2_decap_8
XFILLER_89_7 VPWR VGND sg13g2_fill_2
X_12666_ _06481_ _06479_ VPWR VGND sg13g2_inv_2
X_12597_ _06375_ _06394_ _06412_ _06413_ VPWR VGND sg13g2_a21o_1
X_14405_ _00206_ VGND VPWR _00944_ fpmul.reg_a_out\[2\] clknet_leaf_102_clk sg13g2_dfrbpq_2
X_11617_ VPWR _05522_ _05416_ VGND sg13g2_inv_1
XFILLER_30_389 VPWR VGND sg13g2_decap_4
XFILLER_117_907 VPWR VGND sg13g2_decap_8
X_14336_ _00137_ VGND VPWR _00878_ fpmul.reg_p_out\[0\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_7_541 VPWR VGND sg13g2_fill_1
X_11548_ _05453_ _05438_ fp16_sum_pipe.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_116_417 VPWR VGND sg13g2_fill_2
XFILLER_7_574 VPWR VGND sg13g2_decap_4
XFILLER_116_439 VPWR VGND sg13g2_fill_1
X_11479_ _05392_ fp16_res_pipe.x2\[7\] fpdiv.reg1en.d\[0\] VPWR VGND sg13g2_nand2_1
X_14267_ _00068_ VGND VPWR _00818_ fp16_res_pipe.x2\[0\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_125_984 VPWR VGND sg13g2_decap_8
X_14198_ VPWR _00749_ net105 VGND sg13g2_inv_1
XFILLER_83_1013 VPWR VGND sg13g2_fill_1
XFILLER_83_1002 VPWR VGND sg13g2_decap_8
X_13218_ _06903_ _06899_ _06946_ VPWR VGND sg13g2_nor2_1
X_13149_ _06896_ _06885_ piso.tx_active VPWR VGND sg13g2_nand2_1
XFILLER_44_1008 VPWR VGND sg13g2_decap_4
XFILLER_97_367 VPWR VGND sg13g2_decap_8
XFILLER_97_345 VPWR VGND sg13g2_decap_4
XFILLER_111_166 VPWR VGND sg13g2_decap_8
X_07710_ _02017_ _02006_ acc_sub.exp_mant_logic0.a\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_97_378 VPWR VGND sg13g2_fill_1
XFILLER_78_581 VPWR VGND sg13g2_decap_4
X_08690_ _02905_ _02753_ _02904_ VPWR VGND sg13g2_xnor2_1
XFILLER_78_592 VPWR VGND sg13g2_decap_8
X_07641_ _01954_ net1685 net1793 VPWR VGND sg13g2_nand2_1
XFILLER_93_573 VPWR VGND sg13g2_decap_4
XFILLER_81_702 VPWR VGND sg13g2_fill_1
XFILLER_53_415 VPWR VGND sg13g2_decap_4
X_07572_ VGND VPWR _01806_ _01809_ _01886_ _01805_ sg13g2_a21oi_1
XFILLER_19_692 VPWR VGND sg13g2_fill_2
XFILLER_25_117 VPWR VGND sg13g2_fill_2
XFILLER_25_139 VPWR VGND sg13g2_fill_2
X_09311_ VPWR _03464_ _03402_ VGND sg13g2_inv_1
XFILLER_80_289 VPWR VGND sg13g2_fill_2
XFILLER_80_278 VPWR VGND sg13g2_fill_2
XFILLER_62_982 VPWR VGND sg13g2_fill_2
XFILLER_34_673 VPWR VGND sg13g2_decap_4
X_09242_ _03393_ _03395_ _03396_ VPWR VGND sg13g2_nor2_1
X_09173_ _03338_ VPWR _01289_ VGND net1901 _03337_ sg13g2_o21ai_1
X_08124_ _02261_ _02340_ _02386_ VPWR VGND sg13g2_nor2_1
XFILLER_31_28 VPWR VGND sg13g2_decap_8
XFILLER_119_277 VPWR VGND sg13g2_fill_1
XFILLER_119_266 VPWR VGND sg13g2_decap_8
XFILLER_116_940 VPWR VGND sg13g2_decap_8
XFILLER_107_439 VPWR VGND sg13g2_fill_1
XFILLER_103_9 VPWR VGND sg13g2_fill_1
X_08055_ _02315_ _02320_ _02321_ VPWR VGND sg13g2_nor2_1
XFILLER_122_409 VPWR VGND sg13g2_decap_8
Xplace1741 _02648_ net1741 VPWR VGND sg13g2_buf_2
Xplace1730 _06571_ net1730 VPWR VGND sg13g2_buf_2
Xplace1752 net1751 net1752 VPWR VGND sg13g2_buf_2
Xplace1763 _03988_ net1763 VPWR VGND sg13g2_buf_2
Xplace1785 _01490_ net1785 VPWR VGND sg13g2_buf_2
Xplace1796 acc_sub.reg1en.q\[0\] net1796 VPWR VGND sg13g2_buf_2
XFILLER_89_857 VPWR VGND sg13g2_decap_8
Xplace1774 _02179_ net1774 VPWR VGND sg13g2_buf_2
XFILLER_103_645 VPWR VGND sg13g2_fill_2
XFILLER_102_144 VPWR VGND sg13g2_fill_1
XFILLER_88_345 VPWR VGND sg13g2_decap_4
X_08957_ _03143_ _03142_ acc_sub.add_renorm0.exp\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_102_188 VPWR VGND sg13g2_fill_1
XFILLER_97_890 VPWR VGND sg13g2_decap_8
XFILLER_69_581 VPWR VGND sg13g2_decap_8
XFILLER_57_710 VPWR VGND sg13g2_decap_8
XFILLER_56_14 VPWR VGND sg13g2_decap_8
XFILLER_5_1013 VPWR VGND sg13g2_fill_1
X_08888_ _03062_ _03030_ _03075_ VPWR VGND sg13g2_nor2_1
X_07908_ fp16_sum_pipe.exp_mant_logic0.b\[14\] _02179_ _02183_ VPWR VGND sg13g2_nor2_1
X_07839_ _02132_ _02134_ _02135_ VPWR VGND sg13g2_nor2_1
XFILLER_56_69 VPWR VGND sg13g2_decap_4
XFILLER_29_456 VPWR VGND sg13g2_decap_8
XFILLER_29_467 VPWR VGND sg13g2_decap_8
XFILLER_112_42 VPWR VGND sg13g2_decap_8
XFILLER_44_448 VPWR VGND sg13g2_decap_4
X_10850_ VGND VPWR _04793_ net1825 _04862_ _04861_ sg13g2_a21oi_1
XFILLER_44_459 VPWR VGND sg13g2_fill_2
XFILLER_25_662 VPWR VGND sg13g2_decap_8
XFILLER_72_68 VPWR VGND sg13g2_fill_1
XFILLER_72_57 VPWR VGND sg13g2_fill_2
XFILLER_24_150 VPWR VGND sg13g2_fill_2
X_10781_ _04793_ _03580_ _04778_ VPWR VGND sg13g2_xnor2_1
X_12520_ VGND VPWR _03603_ net1951 _00949_ _06345_ sg13g2_a21oi_1
X_12451_ _06296_ _05876_ fpmul.seg_reg0.q\[14\] VPWR VGND sg13g2_nand2_1
X_11402_ _05346_ net1707 fpdiv.div_out\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_125_203 VPWR VGND sg13g2_decap_8
X_14121_ VPWR _00672_ net99 VGND sg13g2_inv_1
X_12382_ VPWR _06228_ _06227_ VGND sg13g2_inv_1
XFILLER_115_0 VPWR VGND sg13g2_decap_8
XFILLER_67_1008 VPWR VGND sg13g2_decap_4
X_11333_ _01078_ _05286_ _05287_ VPWR VGND sg13g2_nand2_1
XFILLER_4_511 VPWR VGND sg13g2_decap_8
XFILLER_122_910 VPWR VGND sg13g2_decap_8
X_14052_ VPWR _00603_ net87 VGND sg13g2_inv_1
X_11264_ _05226_ _05106_ _05227_ VPWR VGND sg13g2_nor2_2
X_13003_ VGND VPWR net1755 fpmul.seg_reg0.q\[12\] _06771_ _06770_ sg13g2_a21oi_1
X_10215_ _04288_ _04156_ _04289_ VPWR VGND sg13g2_nor2_1
XFILLER_97_76 VPWR VGND sg13g2_decap_4
X_11195_ _05163_ net1808 net1655 _05075_ net1810 VPWR VGND sg13g2_a22oi_1
XFILLER_0_750 VPWR VGND sg13g2_decap_8
XFILLER_122_987 VPWR VGND sg13g2_decap_8
XFILLER_94_315 VPWR VGND sg13g2_decap_8
XFILLER_67_529 VPWR VGND sg13g2_fill_1
X_10146_ _04128_ _04142_ net1662 _04227_ VPWR VGND sg13g2_nand3_1
X_14954_ _00755_ VGND VPWR _01474_ acc_sub.add_renorm0.exp\[6\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_2
X_10077_ _01210_ _04162_ _04163_ VPWR VGND sg13g2_nand2_1
XFILLER_36_927 VPWR VGND sg13g2_decap_8
X_13905_ VPWR _00456_ net8 VGND sg13g2_inv_1
X_14885_ _00686_ VGND VPWR _01405_ acc_sub.exp_mant_logic0.b\[11\] clknet_leaf_54_clk
+ sg13g2_dfrbpq_2
XFILLER_35_437 VPWR VGND sg13g2_fill_2
XFILLER_29_990 VPWR VGND sg13g2_decap_8
XFILLER_63_779 VPWR VGND sg13g2_fill_2
XFILLER_62_256 VPWR VGND sg13g2_fill_1
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_16_640 VPWR VGND sg13g2_fill_2
X_13836_ VPWR _00387_ net14 VGND sg13g2_inv_1
X_13767_ VPWR _00318_ net59 VGND sg13g2_inv_1
X_10979_ fp16_sum_pipe.exp_mant_logic0.b\[15\] fp16_res_pipe.x2\[15\] net1930 _01120_
+ VPWR VGND sg13g2_mux2_1
XFILLER_15_161 VPWR VGND sg13g2_decap_8
X_12718_ _06524_ _06433_ _06437_ VPWR VGND sg13g2_nand2b_1
X_13698_ VPWR _00249_ net54 VGND sg13g2_inv_1
X_12649_ _06417_ _06464_ _06465_ VPWR VGND sg13g2_nor2_1
XFILLER_50_1012 VPWR VGND sg13g2_fill_2
XFILLER_12_890 VPWR VGND sg13g2_decap_8
XFILLER_31_698 VPWR VGND sg13g2_fill_2
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_116_236 VPWR VGND sg13g2_decap_8
X_14319_ _00120_ VGND VPWR _00862_ sipo.word\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_7_393 VPWR VGND sg13g2_fill_1
XFILLER_125_781 VPWR VGND sg13g2_decap_8
XFILLER_113_921 VPWR VGND sg13g2_decap_8
X_09860_ _03969_ net1664 _03845_ VPWR VGND sg13g2_nand2_1
XFILLER_124_280 VPWR VGND sg13g2_decap_8
XFILLER_30_0 VPWR VGND sg13g2_decap_8
X_08811_ _02998_ _02995_ _02997_ VPWR VGND sg13g2_nand2_2
XFILLER_113_998 VPWR VGND sg13g2_decap_8
XFILLER_112_486 VPWR VGND sg13g2_decap_8
X_09791_ _03905_ _03783_ _03904_ VPWR VGND sg13g2_nand2b_1
XFILLER_86_827 VPWR VGND sg13g2_decap_8
XFILLER_100_659 VPWR VGND sg13g2_fill_1
XFILLER_85_359 VPWR VGND sg13g2_decap_4
X_08742_ VPWR _02941_ acc_sum.exp_mant_logic0.a\[11\] VGND sg13g2_inv_1
XFILLER_39_754 VPWR VGND sg13g2_decap_8
X_08673_ _02889_ net1671 _02890_ VPWR VGND sg13g2_nor2_1
XFILLER_66_562 VPWR VGND sg13g2_fill_2
XFILLER_66_551 VPWR VGND sg13g2_decap_8
X_07624_ _01937_ _01921_ _01938_ VPWR VGND sg13g2_nor2_1
XFILLER_26_28 VPWR VGND sg13g2_decap_8
XFILLER_26_426 VPWR VGND sg13g2_decap_8
XFILLER_26_437 VPWR VGND sg13g2_fill_2
XFILLER_35_960 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_4
X_07555_ net1796 _01869_ _01837_ _01870_ VPWR VGND sg13g2_nand3_1
XFILLER_107_1013 VPWR VGND sg13g2_fill_1
X_07486_ acc_sub.exp_mant_logic0.a\[9\] _01808_ _01809_ VPWR VGND sg13g2_nor2_1
XFILLER_42_49 VPWR VGND sg13g2_decap_8
X_09225_ fp16_res_pipe.op_sign_logic0.mantisa_b\[7\] _03378_ _03379_ VPWR VGND sg13g2_nor2_1
XFILLER_21_153 VPWR VGND sg13g2_decap_8
XFILLER_22_687 VPWR VGND sg13g2_decap_4
XFILLER_10_849 VPWR VGND sg13g2_decap_8
XFILLER_22_698 VPWR VGND sg13g2_decap_8
X_09156_ _03327_ acc_sub.x2\[15\] VPWR VGND sg13g2_inv_8
X_09087_ _03271_ _03261_ _03270_ VPWR VGND sg13g2_nand2_1
XFILLER_108_759 VPWR VGND sg13g2_decap_8
X_08107_ _02370_ fp16_sum_pipe.exp_mant_logic0.a\[4\] net1645 _02343_ fp16_sum_pipe.exp_mant_logic0.a\[6\]
+ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_110_clk clknet_5_10__leaf_clk clknet_leaf_110_clk VPWR VGND sg13g2_buf_8
XFILLER_107_258 VPWR VGND sg13g2_decap_8
X_08038_ _02297_ _02300_ _02303_ _02304_ VPWR VGND sg13g2_nor3_1
XFILLER_122_217 VPWR VGND sg13g2_decap_8
XFILLER_115_280 VPWR VGND sg13g2_decap_4
XFILLER_107_42 VPWR VGND sg13g2_decap_4
XFILLER_104_943 VPWR VGND sg13g2_decap_8
X_10000_ _04051_ _04087_ _04088_ VPWR VGND sg13g2_nor2_1
XFILLER_103_464 VPWR VGND sg13g2_decap_8
XFILLER_77_827 VPWR VGND sg13g2_decap_8
XFILLER_49_529 VPWR VGND sg13g2_decap_8
X_09989_ VGND VPWR _04039_ _04007_ _04077_ _04004_ sg13g2_a21oi_1
XFILLER_88_197 VPWR VGND sg13g2_fill_2
XFILLER_67_79 VPWR VGND sg13g2_decap_8
Xclkbuf_5_5__f_clk clknet_4_2_0_clk clknet_5_5__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_91_318 VPWR VGND sg13g2_fill_2
XFILLER_91_307 VPWR VGND sg13g2_decap_8
XFILLER_85_860 VPWR VGND sg13g2_fill_1
XFILLER_57_573 VPWR VGND sg13g2_decap_8
XFILLER_17_404 VPWR VGND sg13g2_decap_8
XFILLER_18_927 VPWR VGND sg13g2_decap_8
XFILLER_123_63 VPWR VGND sg13g2_decap_8
X_11951_ VPWR _05811_ fpmul.seg_reg0.q\[29\] VGND sg13g2_inv_1
X_11882_ _05771_ net1718 _05770_ VPWR VGND sg13g2_nand2_1
XFILLER_83_45 VPWR VGND sg13g2_fill_2
X_14670_ _00471_ VGND VPWR _01198_ fp16_res_pipe.op_sign_logic0.mantisa_b\[7\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_1
X_10902_ _04912_ _04877_ _04875_ VPWR VGND sg13g2_xnor2_1
XFILLER_72_587 VPWR VGND sg13g2_fill_1
XFILLER_60_727 VPWR VGND sg13g2_decap_4
X_13621_ VPWR _00172_ net65 VGND sg13g2_inv_1
X_10833_ _04840_ _04844_ _04845_ VPWR VGND sg13g2_nor2_1
XFILLER_26_982 VPWR VGND sg13g2_decap_8
X_13552_ VPWR _00103_ net88 VGND sg13g2_inv_1
XFILLER_12_120 VPWR VGND sg13g2_fill_1
XFILLER_13_621 VPWR VGND sg13g2_decap_8
XFILLER_13_632 VPWR VGND sg13g2_fill_1
XFILLER_16_83 VPWR VGND sg13g2_fill_2
XFILLER_25_492 VPWR VGND sg13g2_fill_1
X_12503_ VGND VPWR _05357_ net1953 _00956_ _06335_ sg13g2_a21oi_1
XFILLER_13_665 VPWR VGND sg13g2_fill_1
XFILLER_13_676 VPWR VGND sg13g2_decap_8
X_13483_ VPWR _00034_ net23 VGND sg13g2_inv_1
XFILLER_40_484 VPWR VGND sg13g2_fill_2
X_10695_ _04707_ VPWR _04708_ VGND net1771 _04703_ sg13g2_o21ai_1
X_12434_ _06253_ _06263_ _06280_ VPWR VGND sg13g2_nor2_1
XFILLER_8_168 VPWR VGND sg13g2_decap_8
X_12365_ _06211_ _06202_ _06205_ VPWR VGND sg13g2_nand2_1
XFILLER_66_9 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_101_clk clknet_5_15__leaf_clk clknet_leaf_101_clk VPWR VGND sg13g2_buf_8
X_11316_ _05272_ net1812 net1656 acc_sum.exp_mant_logic0.b\[4\] _05124_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_5_864 VPWR VGND sg13g2_decap_8
XFILLER_4_330 VPWR VGND sg13g2_decap_8
X_14104_ VPWR _00655_ net43 VGND sg13g2_inv_1
X_14035_ VPWR _00586_ net106 VGND sg13g2_inv_1
X_12296_ VPWR _06142_ _06124_ VGND sg13g2_inv_1
XFILLER_79_142 VPWR VGND sg13g2_fill_2
X_11247_ net1663 _05210_ _05211_ VPWR VGND sg13g2_nor2b_2
XFILLER_122_784 VPWR VGND sg13g2_decap_8
XFILLER_110_913 VPWR VGND sg13g2_decap_8
XFILLER_67_315 VPWR VGND sg13g2_decap_8
XFILLER_0_591 VPWR VGND sg13g2_decap_8
X_10129_ _04211_ _04210_ net1746 VPWR VGND sg13g2_nand2_1
XFILLER_48_562 VPWR VGND sg13g2_fill_1
XFILLER_48_551 VPWR VGND sg13g2_decap_8
X_14937_ _00738_ VGND VPWR _01457_ acc_sub.exp_mant_logic0.a\[5\] clknet_leaf_56_clk
+ sg13g2_dfrbpq_2
XFILLER_75_381 VPWR VGND sg13g2_fill_1
XFILLER_35_212 VPWR VGND sg13g2_decap_8
XFILLER_36_757 VPWR VGND sg13g2_fill_1
X_14868_ _00669_ VGND VPWR _01392_ fp16_sum_pipe.op_sign_logic0.s_b clknet_leaf_111_clk
+ sg13g2_dfrbpq_1
XFILLER_50_204 VPWR VGND sg13g2_fill_1
X_13819_ VPWR _00370_ net62 VGND sg13g2_inv_1
XFILLER_35_267 VPWR VGND sg13g2_decap_8
XFILLER_17_982 VPWR VGND sg13g2_decap_8
X_07340_ _01701_ _01597_ _01582_ VPWR VGND sg13g2_xnor2_1
X_14799_ _00600_ VGND VPWR _01323_ acc_sum.exp_mant_logic0.a\[12\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_51_749 VPWR VGND sg13g2_decap_8
XFILLER_16_481 VPWR VGND sg13g2_decap_4
XFILLER_32_985 VPWR VGND sg13g2_decap_8
X_09010_ _03196_ _03194_ _03195_ VPWR VGND sg13g2_nand2_1
X_07271_ _01640_ net1783 acc_sub.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_78_0 VPWR VGND sg13g2_decap_8
XFILLER_117_545 VPWR VGND sg13g2_decap_8
XFILLER_117_534 VPWR VGND sg13g2_decap_8
XFILLER_8_691 VPWR VGND sg13g2_decap_8
XFILLER_99_930 VPWR VGND sg13g2_decap_8
X_09912_ _03993_ _03998_ _04003_ _04008_ _04009_ VPWR VGND sg13g2_nor4_1
XFILLER_112_250 VPWR VGND sg13g2_decap_4
XFILLER_101_913 VPWR VGND sg13g2_decap_8
X_09843_ net1769 VPWR _03954_ VGND _03809_ _03953_ sg13g2_o21ai_1
XFILLER_86_602 VPWR VGND sg13g2_decap_8
XFILLER_113_795 VPWR VGND sg13g2_decap_8
X_09774_ _01239_ _03888_ _03889_ VPWR VGND sg13g2_nand2_1
XFILLER_73_307 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
X_08725_ VPWR _02930_ acc_sum.add_renorm0.exp\[1\] VGND sg13g2_inv_1
XFILLER_66_381 VPWR VGND sg13g2_decap_8
XFILLER_54_521 VPWR VGND sg13g2_fill_2
XFILLER_39_595 VPWR VGND sg13g2_decap_8
X_08656_ VGND VPWR _02874_ net1818 _01343_ _02875_ sg13g2_a21oi_1
X_07607_ VPWR _01921_ _01920_ VGND sg13g2_inv_1
X_08587_ VPWR _02810_ _02809_ VGND sg13g2_inv_1
XFILLER_14_407 VPWR VGND sg13g2_decap_4
X_07538_ _01856_ VPWR _01435_ VGND _01804_ _01855_ sg13g2_o21ai_1
XFILLER_41_237 VPWR VGND sg13g2_fill_1
X_07469_ VPWR _01792_ _01791_ VGND sg13g2_inv_1
XFILLER_10_624 VPWR VGND sg13g2_decap_8
XFILLER_23_996 VPWR VGND sg13g2_decap_8
X_09208_ _03363_ fp16_res_pipe.op_sign_logic0.s_a fp16_res_pipe.op_sign_logic0.s_b
+ VPWR VGND sg13g2_xnor2_1
X_10480_ VGND VPWR _04384_ _04526_ _04527_ _04495_ sg13g2_a21oi_1
X_09139_ _03317_ VPWR _03318_ VGND _03070_ _03226_ sg13g2_o21ai_1
XFILLER_6_628 VPWR VGND sg13g2_decap_8
XFILLER_5_105 VPWR VGND sg13g2_decap_8
X_12150_ _05996_ _05994_ _05995_ VPWR VGND sg13g2_nand2_1
XFILLER_118_63 VPWR VGND sg13g2_decap_8
XFILLER_78_23 VPWR VGND sg13g2_fill_1
X_11101_ _05068_ _05069_ _05070_ _05072_ VGND VPWR _05071_ sg13g2_nor4_2
X_12081_ VPWR _05927_ _05926_ VGND sg13g2_inv_1
XFILLER_2_856 VPWR VGND sg13g2_decap_8
XFILLER_104_773 VPWR VGND sg13g2_decap_8
X_11032_ _04998_ _05002_ _05006_ _05010_ _05011_ VPWR VGND sg13g2_nor4_1
XFILLER_1_366 VPWR VGND sg13g2_decap_8
XFILLER_103_294 VPWR VGND sg13g2_decap_8
XFILLER_77_657 VPWR VGND sg13g2_decap_8
XFILLER_49_348 VPWR VGND sg13g2_fill_2
XFILLER_49_337 VPWR VGND sg13g2_decap_8
XFILLER_92_616 VPWR VGND sg13g2_decap_4
XFILLER_58_871 VPWR VGND sg13g2_decap_8
XFILLER_94_77 VPWR VGND sg13g2_decap_8
XFILLER_94_66 VPWR VGND sg13g2_fill_2
XFILLER_73_830 VPWR VGND sg13g2_fill_1
X_12983_ _05873_ _05877_ net1755 _06751_ VPWR VGND sg13g2_nor3_2
X_11934_ _05800_ net1879 fpmul.reg_b_out\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_17_234 VPWR VGND sg13g2_decap_4
X_14722_ _00523_ VGND VPWR _01250_ fp16_res_pipe.exp_mant_logic0.a\[9\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_2
XFILLER_72_373 VPWR VGND sg13g2_fill_2
XFILLER_33_738 VPWR VGND sg13g2_decap_8
X_14653_ _00454_ VGND VPWR _01181_ fp16_res_pipe.exp_mant_logic0.b\[6\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_1
X_13604_ VPWR _00155_ net123 VGND sg13g2_inv_1
XFILLER_60_535 VPWR VGND sg13g2_fill_2
XFILLER_45_598 VPWR VGND sg13g2_decap_8
X_11865_ _05761_ VPWR _01020_ VGND _05760_ _05572_ sg13g2_o21ai_1
XFILLER_33_749 VPWR VGND sg13g2_fill_2
XFILLER_14_930 VPWR VGND sg13g2_decap_8
X_11796_ _05698_ _05496_ _05697_ _05696_ _05491_ VPWR VGND sg13g2_a22oi_1
X_10816_ _04828_ _04826_ _04827_ VPWR VGND sg13g2_nand2_1
X_14584_ _00385_ VGND VPWR _01116_ fp16_sum_pipe.exp_mant_logic0.b\[11\] clknet_leaf_134_clk
+ sg13g2_dfrbpq_1
X_13535_ VPWR _00086_ net85 VGND sg13g2_inv_1
XFILLER_43_70 VPWR VGND sg13g2_decap_8
XFILLER_9_433 VPWR VGND sg13g2_decap_4
XFILLER_13_484 VPWR VGND sg13g2_decap_8
X_10747_ _04759_ VPWR _04760_ VGND fp16_res_pipe.seg_reg1.q\[21\] _04756_ sg13g2_o21ai_1
X_13466_ _07112_ VPWR _00771_ VGND _06939_ net1753 sg13g2_o21ai_1
X_10678_ _04691_ _04689_ _04690_ VPWR VGND sg13g2_xnor2_1
X_12417_ _06263_ _06260_ _06261_ VPWR VGND sg13g2_xnor2_1
XFILLER_127_876 VPWR VGND sg13g2_decap_8
X_13397_ acc_sub.x2\[0\] _07055_ _07075_ VPWR VGND sg13g2_nor2_1
XFILLER_114_537 VPWR VGND sg13g2_fill_1
X_12348_ _06194_ _06191_ _06193_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_672 VPWR VGND sg13g2_decap_8
XFILLER_99_248 VPWR VGND sg13g2_decap_8
X_12279_ _06125_ _06122_ _06123_ VPWR VGND sg13g2_nand2_1
XFILLER_5_694 VPWR VGND sg13g2_fill_1
XFILLER_4_182 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
XFILLER_110_710 VPWR VGND sg13g2_fill_1
X_14018_ VPWR _00569_ net22 VGND sg13g2_inv_1
XFILLER_96_955 VPWR VGND sg13g2_decap_8
XFILLER_95_476 VPWR VGND sg13g2_decap_8
XFILLER_95_465 VPWR VGND sg13g2_decap_8
XFILLER_110_787 VPWR VGND sg13g2_decap_8
XFILLER_67_178 VPWR VGND sg13g2_fill_2
X_08510_ VPWR _02734_ acc_sum.op_sign_logic0.mantisa_b\[7\] VGND sg13g2_inv_1
XFILLER_64_841 VPWR VGND sg13g2_decap_8
X_09490_ _03611_ fp16_res_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_inv_2
X_08441_ _02675_ fpdiv.divider0.divisor_reg\[9\] fpdiv.divider0.remainder_reg\[9\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_91_660 VPWR VGND sg13g2_decap_4
XFILLER_36_587 VPWR VGND sg13g2_decap_8
XFILLER_63_384 VPWR VGND sg13g2_decap_8
X_08372_ VGND VPWR _02610_ _02614_ _02615_ _02591_ sg13g2_a21oi_1
XFILLER_51_579 VPWR VGND sg13g2_decap_8
X_07323_ _01686_ net1666 _01626_ VPWR VGND sg13g2_nand2_1
X_07254_ VGND VPWR _01586_ _01551_ _01624_ _01623_ sg13g2_a21oi_1
XFILLER_118_810 VPWR VGND sg13g2_decap_8
XFILLER_20_955 VPWR VGND sg13g2_decap_8
XFILLER_31_292 VPWR VGND sg13g2_decap_4
X_07185_ acc_sub.op_sign_logic0.mantisa_b\[3\] _01556_ _01557_ VPWR VGND sg13g2_nor2_1
XFILLER_117_331 VPWR VGND sg13g2_fill_1
XFILLER_118_887 VPWR VGND sg13g2_decap_8
XFILLER_2_119 VPWR VGND sg13g2_decap_8
XFILLER_105_559 VPWR VGND sg13g2_decap_8
XFILLER_87_900 VPWR VGND sg13g2_fill_2
XFILLER_101_743 VPWR VGND sg13g2_decap_8
XFILLER_98_270 VPWR VGND sg13g2_fill_2
XFILLER_87_944 VPWR VGND sg13g2_decap_8
X_09826_ _03648_ VPWR _03938_ VGND _03871_ _03937_ sg13g2_o21ai_1
XFILLER_59_679 VPWR VGND sg13g2_fill_1
XFILLER_58_156 VPWR VGND sg13g2_fill_1
X_09757_ _03838_ _03872_ _03873_ VPWR VGND sg13g2_nor2_1
XFILLER_101_798 VPWR VGND sg13g2_fill_2
XFILLER_100_275 VPWR VGND sg13g2_fill_1
XFILLER_58_167 VPWR VGND sg13g2_decap_8
X_08708_ VGND VPWR _02803_ _02918_ _01335_ _02919_ sg13g2_a21oi_1
XFILLER_73_148 VPWR VGND sg13g2_decap_8
XFILLER_55_841 VPWR VGND sg13g2_decap_4
X_09688_ VPWR _03804_ _03803_ VGND sg13g2_inv_1
XFILLER_70_822 VPWR VGND sg13g2_fill_1
XFILLER_70_800 VPWR VGND sg13g2_fill_2
XFILLER_55_896 VPWR VGND sg13g2_fill_1
XFILLER_54_373 VPWR VGND sg13g2_decap_8
XFILLER_42_502 VPWR VGND sg13g2_decap_4
XFILLER_14_204 VPWR VGND sg13g2_decap_8
X_08639_ net1818 acc_sum.add_renorm0.mantisa\[10\] _02861_ VPWR VGND sg13g2_nor2_1
XFILLER_42_524 VPWR VGND sg13g2_decap_8
XFILLER_15_738 VPWR VGND sg13g2_fill_2
XFILLER_120_42 VPWR VGND sg13g2_decap_8
Xfanout30 net31 net30 VPWR VGND sg13g2_buf_2
X_11650_ _05554_ VPWR _05555_ VGND _05498_ _05552_ sg13g2_o21ai_1
XFILLER_80_57 VPWR VGND sg13g2_decap_8
Xfanout74 net76 net74 VPWR VGND sg13g2_buf_2
Xfanout63 net67 net63 VPWR VGND sg13g2_buf_2
Xfanout52 net55 net52 VPWR VGND sg13g2_buf_2
Xfanout41 net42 net41 VPWR VGND sg13g2_buf_1
X_10601_ _04614_ fp16_res_pipe.add_renorm0.mantisa\[11\] fp16_res_pipe.add_renorm0.mantisa\[7\]
+ VPWR VGND sg13g2_nand2_1
X_11581_ _05485_ _05470_ _05435_ _05462_ _05486_ VPWR VGND sg13g2_nor4_1
Xfanout96 net107 net96 VPWR VGND sg13g2_buf_2
Xfanout85 net86 net85 VPWR VGND sg13g2_buf_2
X_10532_ _04572_ _04423_ _04571_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_966 VPWR VGND sg13g2_decap_8
XFILLER_22_281 VPWR VGND sg13g2_fill_2
XFILLER_109_821 VPWR VGND sg13g2_decap_8
XFILLER_7_937 VPWR VGND sg13g2_decap_8
XFILLER_13_84 VPWR VGND sg13g2_decap_8
XFILLER_124_802 VPWR VGND sg13g2_decap_8
XFILLER_108_353 VPWR VGND sg13g2_decap_4
X_13251_ _06973_ _06974_ _06971_ _06975_ VPWR VGND sg13g2_nand3_1
X_10463_ VGND VPWR _04510_ _04436_ _04511_ _04435_ sg13g2_a21oi_1
XFILLER_13_95 VPWR VGND sg13g2_fill_2
XFILLER_123_301 VPWR VGND sg13g2_decap_8
X_12202_ _06042_ _06047_ _06041_ _06048_ VPWR VGND sg13g2_nand3_1
X_13182_ _06922_ VPWR _00865_ VGND _06920_ net1715 sg13g2_o21ai_1
X_10394_ _04437_ _04443_ _04444_ VPWR VGND sg13g2_nor2_1
X_12133_ _05907_ _05931_ _05979_ VPWR VGND sg13g2_nor2_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_124_879 VPWR VGND sg13g2_decap_8
XFILLER_111_518 VPWR VGND sg13g2_fill_2
X_12064_ VGND VPWR _05882_ _05887_ _05910_ _05909_ sg13g2_a21oi_1
XFILLER_2_675 VPWR VGND sg13g2_fill_1
XFILLER_104_570 VPWR VGND sg13g2_decap_4
XFILLER_89_292 VPWR VGND sg13g2_decap_8
XFILLER_77_432 VPWR VGND sg13g2_decap_8
XFILLER_77_421 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_77_454 VPWR VGND sg13g2_decap_8
XFILLER_65_605 VPWR VGND sg13g2_fill_1
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_93_947 VPWR VGND sg13g2_decap_8
XFILLER_65_638 VPWR VGND sg13g2_decap_8
XFILLER_38_70 VPWR VGND sg13g2_decap_8
X_14705_ _00506_ VGND VPWR _01233_ acc_sum.y\[8\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_12966_ _06735_ _06736_ _06726_ _00895_ VPWR VGND sg13g2_nand3_1
XFILLER_61_811 VPWR VGND sg13g2_fill_1
XFILLER_45_351 VPWR VGND sg13g2_decap_8
XFILLER_73_682 VPWR VGND sg13g2_fill_1
X_12897_ acc\[6\] net1907 _03983_ _06673_ VPWR VGND sg13g2_nand3_1
XFILLER_72_170 VPWR VGND sg13g2_fill_1
X_11917_ _05788_ VPWR _00995_ VGND net1881 _05787_ sg13g2_o21ai_1
XFILLER_61_866 VPWR VGND sg13g2_fill_2
X_14636_ _00437_ VGND VPWR _01168_ fp16_sum_pipe.add_renorm0.mantisa\[7\] clknet_leaf_109_clk
+ sg13g2_dfrbpq_2
X_11848_ _05746_ _05491_ _05616_ VPWR VGND sg13g2_nand2_1
XFILLER_33_557 VPWR VGND sg13g2_decap_8
X_14567_ _00368_ VGND VPWR _01103_ acc_sum.op_sign_logic0.s_b clknet_leaf_32_clk sg13g2_dfrbpq_1
XFILLER_14_793 VPWR VGND sg13g2_fill_2
X_13518_ VPWR _00069_ net85 VGND sg13g2_inv_1
X_11779_ _05627_ _05610_ _05642_ _05682_ VPWR VGND sg13g2_nand3_1
X_14498_ _00299_ VGND VPWR _01034_ fpdiv.divider0.divisor\[9\] clknet_leaf_84_clk
+ sg13g2_dfrbpq_1
XFILLER_115_802 VPWR VGND sg13g2_decap_8
Xclkload11 clknet_5_23__leaf_clk clkload11/X VPWR VGND sg13g2_buf_8
Xclkload33 clknet_leaf_3_clk clkload33/X VPWR VGND sg13g2_buf_8
X_13449_ _07104_ net1754 sipo.shift_reg\[9\] VPWR VGND sg13g2_nand2_1
Xclkload22 clkload22/Y clknet_leaf_11_clk VPWR VGND sg13g2_inv_2
Xclkload44 clkload44/Y clknet_leaf_117_clk VPWR VGND sg13g2_inv_8
XFILLER_126_161 VPWR VGND sg13g2_decap_8
XFILLER_114_312 VPWR VGND sg13g2_decap_8
Xclkload77 clknet_leaf_52_clk clkload77/Y VPWR VGND sg13g2_inv_4
Xclkload66 clkload66/Y clknet_leaf_102_clk VPWR VGND sg13g2_inv_8
Xclkload55 clkload55/Y clknet_leaf_96_clk VPWR VGND sg13g2_inv_2
Xclkload88 VPWR clkload88/Y clknet_leaf_42_clk VGND sg13g2_inv_1
Xclkload99 VPWR clkload99/Y clknet_leaf_80_clk VGND sg13g2_inv_1
X_08990_ _03176_ _03175_ _03086_ VPWR VGND sg13g2_xnor2_1
XFILLER_115_879 VPWR VGND sg13g2_decap_8
XFILLER_114_367 VPWR VGND sg13g2_decap_8
XFILLER_123_890 VPWR VGND sg13g2_decap_8
X_07941_ _02216_ fp16_sum_pipe.exp_mant_logic0.b\[7\] VPWR VGND sg13g2_inv_2
XFILLER_110_540 VPWR VGND sg13g2_fill_1
XFILLER_95_240 VPWR VGND sg13g2_fill_2
X_07872_ _02163_ net1888 acc_sub.x2\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_69_977 VPWR VGND sg13g2_decap_8
XFILLER_110_573 VPWR VGND sg13g2_decap_8
X_09611_ _03728_ _03727_ _03707_ VPWR VGND sg13g2_nand2b_1
XFILLER_56_627 VPWR VGND sg13g2_decap_4
X_09542_ _03635_ _03658_ _03659_ VPWR VGND sg13g2_nor2_1
XFILLER_110_595 VPWR VGND sg13g2_fill_2
XFILLER_37_841 VPWR VGND sg13g2_decap_8
XFILLER_70_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_90_clk clknet_5_24__leaf_clk clknet_leaf_90_clk VPWR VGND sg13g2_buf_8
XFILLER_37_896 VPWR VGND sg13g2_decap_8
X_09473_ _03600_ acc_sub.x2\[9\] net1912 VPWR VGND sg13g2_nand2_1
XFILLER_34_28 VPWR VGND sg13g2_decap_8
XFILLER_24_513 VPWR VGND sg13g2_fill_2
XFILLER_24_546 VPWR VGND sg13g2_decap_8
X_08424_ VPWR _02658_ fpdiv.divider0.remainder_reg\[7\] VGND sg13g2_inv_1
XFILLER_51_332 VPWR VGND sg13g2_decap_8
X_08355_ _02598_ _02596_ _02597_ VPWR VGND sg13g2_nand2_2
X_07306_ _01542_ _01571_ _01671_ VPWR VGND sg13g2_nor2_1
XFILLER_20_741 VPWR VGND sg13g2_decap_8
Xclkload5 clknet_5_11__leaf_clk clkload5/X VPWR VGND sg13g2_buf_8
XFILLER_109_128 VPWR VGND sg13g2_decap_8
XFILLER_109_106 VPWR VGND sg13g2_decap_8
XFILLER_50_49 VPWR VGND sg13g2_decap_8
X_08286_ _02534_ fp16_sum_pipe.exp_mant_logic0.b\[6\] _02408_ _02472_ _02332_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_20_763 VPWR VGND sg13g2_fill_2
X_07237_ _01608_ _01607_ _01528_ VPWR VGND sg13g2_nand2_1
XFILLER_119_7 VPWR VGND sg13g2_decap_8
X_07168_ acc_sub.op_sign_logic0.mantisa_a\[4\] _01539_ _01540_ VPWR VGND sg13g2_nor2_1
XFILLER_117_161 VPWR VGND sg13g2_decap_8
XFILLER_3_406 VPWR VGND sg13g2_decap_8
Xclkbuf_5_30__f_clk clknet_4_15_0_clk clknet_5_30__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_121_805 VPWR VGND sg13g2_decap_8
XFILLER_79_719 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_120_315 VPWR VGND sg13g2_fill_1
XFILLER_87_730 VPWR VGND sg13g2_decap_8
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
XFILLER_115_42 VPWR VGND sg13g2_decap_8
XFILLER_101_540 VPWR VGND sg13g2_decap_8
XFILLER_75_903 VPWR VGND sg13g2_fill_1
XFILLER_59_432 VPWR VGND sg13g2_fill_1
X_09809_ _03908_ _03907_ _03922_ VPWR VGND sg13g2_nor2_1
XFILLER_75_35 VPWR VGND sg13g2_decap_8
XFILLER_59_498 VPWR VGND sg13g2_decap_8
XFILLER_19_307 VPWR VGND sg13g2_fill_2
XFILLER_101_595 VPWR VGND sg13g2_decap_8
X_12820_ _06603_ net1716 _00018_ VPWR VGND sg13g2_nand2_1
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_90_939 VPWR VGND sg13g2_decap_8
XFILLER_55_660 VPWR VGND sg13g2_fill_2
XFILLER_43_800 VPWR VGND sg13g2_fill_2
X_12751_ _06543_ fp16_res_pipe.x2\[6\] net1955 VPWR VGND sg13g2_nand2_1
XFILLER_42_310 VPWR VGND sg13g2_fill_2
XFILLER_15_524 VPWR VGND sg13g2_fill_2
XFILLER_15_535 VPWR VGND sg13g2_decap_8
XFILLER_28_896 VPWR VGND sg13g2_decap_8
X_12682_ VGND VPWR _06464_ _06493_ _06494_ net1735 sg13g2_a21oi_1
XFILLER_70_641 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_81_clk clknet_5_26__leaf_clk clknet_leaf_81_clk VPWR VGND sg13g2_buf_8
XFILLER_43_888 VPWR VGND sg13g2_fill_1
XFILLER_42_332 VPWR VGND sg13g2_decap_8
X_11702_ _05606_ fp16_sum_pipe.add_renorm0.exp\[5\] _05578_ VPWR VGND sg13g2_xnor2_1
XFILLER_15_546 VPWR VGND sg13g2_fill_2
XFILLER_15_579 VPWR VGND sg13g2_decap_8
X_14421_ _00222_ VGND VPWR _00960_ fpmul.seg_reg0.q\[6\] clknet_leaf_78_clk sg13g2_dfrbpq_1
XFILLER_43_899 VPWR VGND sg13g2_fill_2
XFILLER_42_398 VPWR VGND sg13g2_fill_1
X_11633_ _05538_ _05412_ _05526_ VPWR VGND sg13g2_nand2_1
X_14352_ _00153_ VGND VPWR _00894_ _00005_ clknet_leaf_82_clk sg13g2_dfrbpq_1
X_11564_ VPWR _05469_ _05468_ VGND sg13g2_inv_1
X_13303_ _07014_ _06952_ _07015_ VPWR VGND sg13g2_nor2_1
X_14283_ _00084_ VGND VPWR _07116_ fpmul.reg1en.d\[0\] clknet_leaf_53_clk sg13g2_dfrbpq_2
XFILLER_7_767 VPWR VGND sg13g2_decap_8
XFILLER_6_233 VPWR VGND sg13g2_decap_8
X_10515_ _04557_ net1673 _04431_ VPWR VGND sg13g2_nand2_1
X_11495_ _05399_ VPWR _05400_ VGND net1841 _05398_ sg13g2_o21ai_1
X_13234_ _02592_ VPWR _06959_ VGND _02598_ _06958_ sg13g2_o21ai_1
X_10446_ _04494_ VPWR _04495_ VGND _04453_ _04493_ sg13g2_o21ai_1
XFILLER_124_665 VPWR VGND sg13g2_decap_8
X_13165_ _06910_ VPWR _00870_ VGND _06902_ _06906_ sg13g2_o21ai_1
XFILLER_3_973 VPWR VGND sg13g2_decap_8
X_10377_ VPWR _04427_ _04426_ VGND sg13g2_inv_1
XFILLER_123_175 VPWR VGND sg13g2_decap_8
XFILLER_112_838 VPWR VGND sg13g2_decap_8
X_13096_ VPWR _06856_ _06801_ VGND sg13g2_inv_1
XFILLER_69_218 VPWR VGND sg13g2_decap_8
X_12116_ net1858 net1860 _05952_ _05962_ VPWR VGND fpmul.reg_b_out\[5\] sg13g2_nand4_1
XFILLER_34_7 VPWR VGND sg13g2_decap_8
XFILLER_2_472 VPWR VGND sg13g2_decap_8
XFILLER_78_763 VPWR VGND sg13g2_decap_8
X_12047_ _05893_ net1858 fpmul.reg_b_out\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_93_711 VPWR VGND sg13g2_fill_1
XFILLER_66_947 VPWR VGND sg13g2_decap_8
XFILLER_66_925 VPWR VGND sg13g2_decap_8
XFILLER_65_413 VPWR VGND sg13g2_fill_2
XFILLER_65_402 VPWR VGND sg13g2_decap_8
XFILLER_38_638 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_77_284 VPWR VGND sg13g2_fill_1
XFILLER_37_126 VPWR VGND sg13g2_fill_2
XFILLER_92_276 VPWR VGND sg13g2_decap_4
XFILLER_92_243 VPWR VGND sg13g2_fill_2
XFILLER_80_405 VPWR VGND sg13g2_decap_4
XFILLER_53_608 VPWR VGND sg13g2_fill_1
XFILLER_37_159 VPWR VGND sg13g2_fill_1
X_13998_ VPWR _00549_ net9 VGND sg13g2_inv_1
XFILLER_1_98 VPWR VGND sg13g2_decap_8
X_12949_ VPWR _06721_ fpmul.reg_p_out\[2\] VGND sg13g2_inv_1
XFILLER_34_822 VPWR VGND sg13g2_fill_1
XFILLER_33_310 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_72_clk clknet_5_30__leaf_clk clknet_leaf_72_clk VPWR VGND sg13g2_buf_8
XFILLER_60_140 VPWR VGND sg13g2_fill_1
XFILLER_34_866 VPWR VGND sg13g2_decap_8
X_14619_ _00420_ VGND VPWR _01151_ fp16_sum_pipe.exp_mant_logic0.a\[14\] clknet_leaf_134_clk
+ sg13g2_dfrbpq_2
X_08140_ _02401_ fp16_sum_pipe.exp_mant_logic0.a\[5\] net1658 fp16_sum_pipe.exp_mant_logic0.a\[3\]
+ net1659 VPWR VGND sg13g2_a22oi_1
XFILLER_33_398 VPWR VGND sg13g2_fill_1
XFILLER_119_415 VPWR VGND sg13g2_decap_8
Xclkload111 clkload111/Y clknet_leaf_74_clk VPWR VGND sg13g2_inv_2
Xclkload100 clknet_leaf_83_clk clkload100/Y VPWR VGND sg13g2_inv_4
X_08071_ _02336_ _02315_ _02337_ VPWR VGND sg13g2_nor2_1
XFILLER_115_610 VPWR VGND sg13g2_fill_1
XFILLER_106_109 VPWR VGND sg13g2_fill_1
Xplace1901 net1900 net1901 VPWR VGND sg13g2_buf_2
XFILLER_60_0 VPWR VGND sg13g2_fill_2
Xplace1912 net1911 net1912 VPWR VGND sg13g2_buf_2
XFILLER_127_492 VPWR VGND sg13g2_decap_8
Xplace1945 net1944 net1945 VPWR VGND sg13g2_buf_2
Xplace1923 net1922 net1923 VPWR VGND sg13g2_buf_2
Xplace1934 net1933 net1934 VPWR VGND sg13g2_buf_2
XFILLER_115_665 VPWR VGND sg13g2_decap_8
Xplace1956 net1954 net1956 VPWR VGND sg13g2_buf_2
X_08973_ _03159_ _03146_ acc_sub.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_114_186 VPWR VGND sg13g2_decap_8
XFILLER_114_175 VPWR VGND sg13g2_decap_8
XFILLER_69_752 VPWR VGND sg13g2_decap_8
XFILLER_57_903 VPWR VGND sg13g2_fill_2
X_07924_ fp16_sum_pipe.exp_mant_logic0.b\[12\] _02199_ VPWR VGND sg13g2_inv_4
XFILLER_29_28 VPWR VGND sg13g2_decap_8
XFILLER_84_722 VPWR VGND sg13g2_decap_8
XFILLER_69_785 VPWR VGND sg13g2_decap_8
XFILLER_56_413 VPWR VGND sg13g2_decap_8
X_07855_ _01411_ _02148_ _02149_ VPWR VGND sg13g2_nand2_1
XFILLER_56_435 VPWR VGND sg13g2_fill_2
XFILLER_28_126 VPWR VGND sg13g2_decap_8
X_07786_ _02086_ acc_sub.exp_mant_logic0.b\[3\] net1669 acc_sub.op_sign_logic0.mantisa_b\[6\]
+ net1781 VPWR VGND sg13g2_a22oi_1
XFILLER_25_800 VPWR VGND sg13g2_fill_2
X_09525_ VPWR _03642_ _03627_ VGND sg13g2_inv_1
XFILLER_45_49 VPWR VGND sg13g2_decap_8
XFILLER_36_170 VPWR VGND sg13g2_decap_8
XFILLER_25_822 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_63_clk clknet_5_29__leaf_clk clknet_leaf_63_clk VPWR VGND sg13g2_buf_8
XFILLER_80_972 VPWR VGND sg13g2_decap_8
XFILLER_80_961 VPWR VGND sg13g2_decap_8
X_09456_ VGND VPWR _03327_ net1911 _01256_ _03588_ sg13g2_a21oi_1
XFILLER_25_855 VPWR VGND sg13g2_fill_2
XFILLER_25_866 VPWR VGND sg13g2_fill_1
X_08407_ _02642_ VPWR _01358_ VGND _02589_ _02641_ sg13g2_o21ai_1
XFILLER_52_685 VPWR VGND sg13g2_decap_4
XFILLER_51_173 VPWR VGND sg13g2_fill_1
X_09387_ _03532_ _03534_ _03531_ _01271_ VPWR VGND sg13g2_nand3_1
X_08338_ sipo.word\[10\] sipo.word\[9\] sipo.word\[11\] _02583_ VPWR VGND sipo.word\[8\]
+ sg13g2_nand4_1
X_08269_ _02517_ VPWR _02518_ VGND _02460_ _02322_ sg13g2_o21ai_1
XFILLER_125_429 VPWR VGND sg13g2_fill_2
XFILLER_119_982 VPWR VGND sg13g2_decap_8
X_11280_ _01085_ _05240_ _05241_ VPWR VGND sg13g2_nand2_1
X_10300_ _04368_ net1763 fp16_res_pipe.op_sign_logic0.mantisa_b\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_106_643 VPWR VGND sg13g2_decap_8
XFILLER_3_203 VPWR VGND sg13g2_decap_8
X_10231_ _04299_ _04301_ _04303_ _04304_ VPWR VGND sg13g2_nor3_1
XFILLER_121_602 VPWR VGND sg13g2_decap_8
XFILLER_106_654 VPWR VGND sg13g2_fill_2
XFILLER_10_63 VPWR VGND sg13g2_decap_8
XFILLER_126_63 VPWR VGND sg13g2_decap_8
XFILLER_121_635 VPWR VGND sg13g2_decap_8
XFILLER_120_112 VPWR VGND sg13g2_decap_8
X_10162_ _01204_ _04241_ _04242_ VPWR VGND sg13g2_nand2_1
XFILLER_0_954 VPWR VGND sg13g2_decap_8
X_10093_ _04178_ _04177_ net1746 VPWR VGND sg13g2_nand2_1
XFILLER_120_189 VPWR VGND sg13g2_decap_8
XFILLER_102_871 VPWR VGND sg13g2_decap_8
XFILLER_59_262 VPWR VGND sg13g2_decap_8
XFILLER_47_402 VPWR VGND sg13g2_decap_8
X_13921_ VPWR _00472_ net11 VGND sg13g2_inv_1
X_13852_ VPWR _00403_ net30 VGND sg13g2_inv_1
XFILLER_35_619 VPWR VGND sg13g2_fill_2
X_13783_ VPWR _00334_ net125 VGND sg13g2_inv_1
X_12803_ _06587_ _06586_ net1958 VPWR VGND sg13g2_nand2_1
XFILLER_62_416 VPWR VGND sg13g2_decap_8
X_12734_ _06537_ _06442_ _06428_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_54_clk clknet_5_25__leaf_clk clknet_leaf_54_clk VPWR VGND sg13g2_buf_8
X_10995_ _04983_ VPWR _01112_ VGND net1933 _02216_ sg13g2_o21ai_1
XFILLER_15_321 VPWR VGND sg13g2_decap_8
XFILLER_27_192 VPWR VGND sg13g2_decap_4
XFILLER_42_140 VPWR VGND sg13g2_decap_8
X_12665_ _06480_ VPWR _00940_ VGND _06371_ net1741 sg13g2_o21ai_1
XFILLER_31_858 VPWR VGND sg13g2_decap_8
X_12596_ _06374_ _06373_ _06412_ VPWR VGND sg13g2_and2_1
X_14404_ _00205_ VGND VPWR _00943_ fpmul.reg_a_out\[1\] clknet_leaf_102_clk sg13g2_dfrbpq_1
X_11616_ _05412_ _05520_ _05521_ VPWR VGND sg13g2_nor2_1
XFILLER_30_379 VPWR VGND sg13g2_fill_2
X_14335_ _00136_ VGND VPWR _00877_ piso.tx_bit_counter\[4\] clknet_leaf_57_clk sg13g2_dfrbpq_1
XFILLER_51_81 VPWR VGND sg13g2_decap_8
XFILLER_51_70 VPWR VGND sg13g2_fill_1
X_11547_ _05445_ VPWR _05452_ VGND _05451_ _05409_ sg13g2_o21ai_1
X_14266_ _00067_ VGND VPWR _00817_ acc_sub.x2\[15\] clknet_leaf_50_clk sg13g2_dfrbpq_2
X_11478_ VPWR _05391_ fpdiv.reg_b_out\[7\] VGND sg13g2_inv_1
XFILLER_125_963 VPWR VGND sg13g2_decap_8
XFILLER_124_451 VPWR VGND sg13g2_fill_1
XFILLER_98_814 VPWR VGND sg13g2_fill_2
X_14197_ VPWR _00748_ net90 VGND sg13g2_inv_1
X_13217_ VPWR _06945_ _06898_ VGND sg13g2_inv_1
X_10429_ VPWR _04478_ _04423_ VGND sg13g2_inv_1
XFILLER_98_858 VPWR VGND sg13g2_fill_2
XFILLER_98_847 VPWR VGND sg13g2_decap_8
X_13148_ _06895_ VPWR _00872_ VGND _00005_ _06566_ sg13g2_o21ai_1
XFILLER_3_770 VPWR VGND sg13g2_decap_8
XFILLER_39_903 VPWR VGND sg13g2_decap_8
XFILLER_100_819 VPWR VGND sg13g2_decap_8
X_13079_ _06844_ VPWR _00890_ VGND net1861 _06610_ sg13g2_o21ai_1
XFILLER_120_690 VPWR VGND sg13g2_decap_4
X_07640_ _01953_ _01923_ net1792 VPWR VGND sg13g2_nand2_1
XFILLER_93_552 VPWR VGND sg13g2_decap_8
XFILLER_66_788 VPWR VGND sg13g2_decap_4
XFILLER_26_619 VPWR VGND sg13g2_decap_8
X_07571_ _01811_ _01884_ _01885_ VPWR VGND sg13g2_nor2_1
XFILLER_80_224 VPWR VGND sg13g2_fill_2
XFILLER_66_799 VPWR VGND sg13g2_fill_2
XFILLER_53_438 VPWR VGND sg13g2_decap_8
XFILLER_19_671 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_45_clk clknet_5_22__leaf_clk clknet_leaf_45_clk VPWR VGND sg13g2_buf_8
XFILLER_80_257 VPWR VGND sg13g2_decap_8
XFILLER_53_449 VPWR VGND sg13g2_decap_8
XFILLER_34_652 VPWR VGND sg13g2_decap_8
X_09310_ _03462_ VPWR _03463_ VGND _03405_ _03403_ sg13g2_o21ai_1
XFILLER_34_696 VPWR VGND sg13g2_fill_1
XFILLER_33_140 VPWR VGND sg13g2_decap_8
X_09241_ fp16_res_pipe.op_sign_logic0.mantisa_b\[5\] _03394_ _03395_ VPWR VGND sg13g2_nor2_1
X_09172_ _03338_ acc_sub.x2\[10\] net1900 VPWR VGND sg13g2_nand2_1
XFILLER_119_245 VPWR VGND sg13g2_decap_8
X_08123_ _02269_ _02223_ _02385_ VPWR VGND sg13g2_nor2_1
X_08054_ _02320_ _02319_ _02318_ VPWR VGND sg13g2_nand2b_1
Xplace1720 _07076_ net1720 VPWR VGND sg13g2_buf_2
Xplace1742 _02569_ net1742 VPWR VGND sg13g2_buf_2
Xplace1731 net1730 net1731 VPWR VGND sg13g2_buf_2
Xplace1753 net1752 net1753 VPWR VGND sg13g2_buf_2
XFILLER_116_996 VPWR VGND sg13g2_decap_8
XFILLER_115_462 VPWR VGND sg13g2_fill_1
Xplace1786 net1785 net1786 VPWR VGND sg13g2_buf_2
Xplace1797 acc_sub.reg2en.q\[0\] net1797 VPWR VGND sg13g2_buf_2
XFILLER_102_101 VPWR VGND sg13g2_fill_2
XFILLER_89_836 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_fill_2
XFILLER_1_729 VPWR VGND sg13g2_fill_2
Xplace1764 net1763 net1764 VPWR VGND sg13g2_buf_2
Xplace1775 net1774 net1775 VPWR VGND sg13g2_buf_2
XFILLER_103_668 VPWR VGND sg13g2_decap_4
XFILLER_0_239 VPWR VGND sg13g2_decap_8
X_08956_ _01713_ _03141_ _03142_ VPWR VGND sg13g2_nor2_1
XFILLER_97_880 VPWR VGND sg13g2_decap_4
X_08887_ _03074_ _03071_ _03073_ _03055_ _03001_ VPWR VGND sg13g2_a22oi_1
X_07907_ VPWR _02182_ fp16_sum_pipe.seg_reg0.q\[29\] VGND sg13g2_inv_1
X_07838_ _02133_ VPWR _02134_ VGND _02089_ _02024_ sg13g2_o21ai_1
XFILLER_72_714 VPWR VGND sg13g2_decap_8
XFILLER_112_21 VPWR VGND sg13g2_decap_8
XFILLER_38_980 VPWR VGND sg13g2_decap_8
X_07769_ _02071_ net1640 _02070_ VPWR VGND sg13g2_nand2_1
X_09508_ acc_sum.add_renorm0.mantisa\[8\] acc_sum.add_renorm0.mantisa\[7\] _03624_
+ _03625_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_36_clk clknet_5_21__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_71_235 VPWR VGND sg13g2_decap_4
XFILLER_60_909 VPWR VGND sg13g2_decap_8
XFILLER_25_630 VPWR VGND sg13g2_fill_2
XFILLER_25_641 VPWR VGND sg13g2_fill_2
XFILLER_112_98 VPWR VGND sg13g2_decap_8
XFILLER_71_279 VPWR VGND sg13g2_decap_8
XFILLER_12_302 VPWR VGND sg13g2_fill_2
XFILLER_13_825 VPWR VGND sg13g2_fill_1
XFILLER_12_324 VPWR VGND sg13g2_decap_4
X_09439_ VPWR _03578_ fp16_res_pipe.add_renorm0.exp\[5\] VGND sg13g2_inv_1
X_12450_ net1870 _06289_ _06295_ VPWR VGND _06294_ sg13g2_nand3b_1
XFILLER_8_317 VPWR VGND sg13g2_decap_4
XFILLER_12_346 VPWR VGND sg13g2_decap_8
X_11401_ VPWR _05345_ fpdiv.div_out\[5\] VGND sg13g2_inv_1
X_14120_ VPWR _00671_ net101 VGND sg13g2_inv_1
X_12381_ _06227_ net1859 fpmul.reg_b_out\[1\] VPWR VGND sg13g2_nand2_1
X_11332_ _05287_ acc_sum.exp_mant_logic0.b\[2\] net1681 acc_sum.op_sign_logic0.mantisa_b\[5\]
+ net1762 VPWR VGND sg13g2_a22oi_1
XFILLER_125_259 VPWR VGND sg13g2_decap_8
XFILLER_108_0 VPWR VGND sg13g2_decap_8
X_11263_ _05116_ _05020_ _05119_ _05226_ VPWR VGND _05023_ sg13g2_nand4_1
X_14051_ VPWR _00602_ net22 VGND sg13g2_inv_1
XFILLER_21_95 VPWR VGND sg13g2_decap_4
XFILLER_121_410 VPWR VGND sg13g2_decap_8
XFILLER_107_985 VPWR VGND sg13g2_decap_8
XFILLER_106_462 VPWR VGND sg13g2_decap_8
XFILLER_79_313 VPWR VGND sg13g2_decap_8
X_11194_ _05162_ net1809 _05161_ _05141_ _05073_ VPWR VGND sg13g2_a22oi_1
X_13002_ VPWR _06770_ _06769_ VGND sg13g2_inv_1
X_10214_ _04288_ fp16_res_pipe.exp_mant_logic0.b\[5\] VPWR VGND sg13g2_inv_2
XFILLER_122_966 VPWR VGND sg13g2_decap_8
XFILLER_121_421 VPWR VGND sg13g2_fill_2
XFILLER_79_357 VPWR VGND sg13g2_decap_4
X_10145_ _04225_ VPWR _04226_ VGND _03605_ _04222_ sg13g2_o21ai_1
XFILLER_48_711 VPWR VGND sg13g2_fill_1
X_14953_ _00754_ VGND VPWR _01473_ acc_sub.add_renorm0.exp\[5\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_94_349 VPWR VGND sg13g2_decap_8
X_10076_ _04163_ net1828 net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[8\] net1764
+ VPWR VGND sg13g2_a22oi_1
X_14884_ _00685_ VGND VPWR _01404_ acc_sub.exp_mant_logic0.b\[10\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_2
XFILLER_36_906 VPWR VGND sg13g2_decap_8
X_13904_ VPWR _00455_ net12 VGND sg13g2_inv_1
XFILLER_62_224 VPWR VGND sg13g2_fill_1
XFILLER_46_70 VPWR VGND sg13g2_decap_8
X_13835_ VPWR _00386_ net51 VGND sg13g2_inv_1
Xclkbuf_leaf_27_clk clknet_5_16__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
X_13766_ VPWR _00317_ net115 VGND sg13g2_inv_1
XFILLER_62_268 VPWR VGND sg13g2_fill_2
XFILLER_44_994 VPWR VGND sg13g2_decap_8
X_10978_ _04975_ VPWR _01121_ VGND _04772_ _04759_ sg13g2_o21ai_1
X_12717_ _06521_ _06522_ _06452_ _06523_ VPWR VGND _06425_ sg13g2_nand4_1
X_13697_ VPWR _00248_ net54 VGND sg13g2_inv_1
X_12648_ VPWR _06464_ _06463_ VGND sg13g2_inv_1
XFILLER_62_80 VPWR VGND sg13g2_decap_8
XFILLER_30_165 VPWR VGND sg13g2_decap_8
X_12579_ _06395_ _06375_ _06394_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_11_1008 VPWR VGND sg13g2_decap_4
XFILLER_30_198 VPWR VGND sg13g2_decap_4
XFILLER_116_215 VPWR VGND sg13g2_decap_8
X_14318_ _00119_ VGND VPWR _00861_ sipo.word\[6\] clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_8_895 VPWR VGND sg13g2_decap_8
XFILLER_125_760 VPWR VGND sg13g2_decap_8
XFILLER_113_900 VPWR VGND sg13g2_decap_8
X_14249_ _00050_ VGND VPWR _00800_ instr\[14\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_112_410 VPWR VGND sg13g2_fill_2
X_08810_ _02997_ _02996_ VPWR VGND sg13g2_inv_2
XFILLER_113_977 VPWR VGND sg13g2_decap_8
XFILLER_112_465 VPWR VGND sg13g2_decap_8
X_09790_ VGND VPWR _03902_ _03903_ _03904_ net1803 sg13g2_a21oi_1
XFILLER_98_688 VPWR VGND sg13g2_decap_4
XFILLER_97_176 VPWR VGND sg13g2_fill_1
XFILLER_23_0 VPWR VGND sg13g2_decap_8
X_08741_ _02940_ VPWR _01323_ VGND net1904 _02939_ sg13g2_o21ai_1
X_08672_ VGND VPWR _02769_ _02774_ _02889_ _02771_ sg13g2_a21oi_1
X_07623_ VPWR _01937_ _01936_ VGND sg13g2_inv_1
XFILLER_81_522 VPWR VGND sg13g2_decap_8
XFILLER_66_596 VPWR VGND sg13g2_decap_8
XFILLER_38_276 VPWR VGND sg13g2_decap_8
XFILLER_38_265 VPWR VGND sg13g2_fill_1
XFILLER_27_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_18_clk clknet_5_7__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_19_490 VPWR VGND sg13g2_fill_1
X_07554_ _01868_ _01869_ VPWR VGND sg13g2_inv_4
XFILLER_53_268 VPWR VGND sg13g2_decap_4
XFILLER_41_408 VPWR VGND sg13g2_fill_1
X_07485_ VPWR _01808_ acc_sub.exp_mant_logic0.b\[9\] VGND sg13g2_inv_1
XFILLER_22_633 VPWR VGND sg13g2_decap_8
XFILLER_22_644 VPWR VGND sg13g2_fill_1
XFILLER_42_28 VPWR VGND sg13g2_decap_8
X_09224_ VPWR _03378_ fp16_res_pipe.op_sign_logic0.mantisa_a\[7\] VGND sg13g2_inv_1
XFILLER_10_828 VPWR VGND sg13g2_decap_8
XFILLER_21_187 VPWR VGND sg13g2_decap_8
X_09155_ _03326_ VPWR _01295_ VGND net1773 _03074_ sg13g2_o21ai_1
XFILLER_21_198 VPWR VGND sg13g2_fill_2
X_09086_ _03270_ _03264_ _03269_ VPWR VGND sg13g2_nand2_1
XFILLER_108_738 VPWR VGND sg13g2_decap_8
XFILLER_107_237 VPWR VGND sg13g2_decap_8
X_08106_ _01380_ _02367_ _02369_ VPWR VGND sg13g2_nand2_1
XFILLER_101_7 VPWR VGND sg13g2_fill_2
X_08037_ _02302_ _02190_ _02303_ VPWR VGND sg13g2_xor2_1
XFILLER_116_793 VPWR VGND sg13g2_decap_8
XFILLER_104_922 VPWR VGND sg13g2_decap_8
XFILLER_89_622 VPWR VGND sg13g2_decap_8
XFILLER_89_600 VPWR VGND sg13g2_fill_1
XFILLER_103_443 VPWR VGND sg13g2_decap_8
XFILLER_88_132 VPWR VGND sg13g2_fill_2
XFILLER_88_121 VPWR VGND sg13g2_decap_8
XFILLER_77_806 VPWR VGND sg13g2_fill_2
XFILLER_114_1007 VPWR VGND sg13g2_decap_8
XFILLER_107_98 VPWR VGND sg13g2_decap_8
XFILLER_104_999 VPWR VGND sg13g2_decap_8
XFILLER_103_476 VPWR VGND sg13g2_decap_8
X_09988_ VPWR _04076_ net1703 VGND sg13g2_inv_1
X_08939_ _03126_ _03014_ _03001_ VPWR VGND sg13g2_nand2_1
XFILLER_67_69 VPWR VGND sg13g2_fill_2
XFILLER_123_42 VPWR VGND sg13g2_decap_8
X_11950_ _05810_ VPWR _00984_ VGND net1884 _05809_ sg13g2_o21ai_1
XFILLER_18_906 VPWR VGND sg13g2_decap_8
XFILLER_29_254 VPWR VGND sg13g2_decap_8
X_10901_ _04911_ _04905_ _04910_ VPWR VGND sg13g2_nand2_1
X_11881_ _05770_ _02644_ _05769_ VPWR VGND sg13g2_xnor2_1
XFILLER_45_769 VPWR VGND sg13g2_decap_8
XFILLER_83_79 VPWR VGND sg13g2_decap_4
X_13620_ VPWR _00171_ net66 VGND sg13g2_inv_1
XFILLER_13_600 VPWR VGND sg13g2_decap_8
X_10832_ _04842_ _04843_ _04844_ VPWR VGND sg13g2_nor2_1
XFILLER_26_961 VPWR VGND sg13g2_decap_8
X_13551_ VPWR _00102_ net87 VGND sg13g2_inv_1
XFILLER_41_942 VPWR VGND sg13g2_decap_8
X_10763_ _04653_ _04652_ _04775_ VPWR VGND sg13g2_nor2_2
X_12502_ fpmul.reg_a_out\[14\] net1953 _06335_ VPWR VGND sg13g2_nor2_1
XFILLER_41_986 VPWR VGND sg13g2_decap_8
X_13482_ VPWR _00033_ net23 VGND sg13g2_inv_1
XFILLER_9_648 VPWR VGND sg13g2_fill_2
X_10694_ _03359_ _04706_ _04707_ VPWR VGND _04705_ sg13g2_nand3b_1
XFILLER_126_502 VPWR VGND sg13g2_fill_2
X_12433_ _06279_ _06252_ _06278_ VPWR VGND sg13g2_nand2_1
XFILLER_8_147 VPWR VGND sg13g2_decap_8
X_12364_ _06210_ _06185_ _06209_ VPWR VGND sg13g2_nand2_1
XFILLER_114_719 VPWR VGND sg13g2_decap_4
X_11315_ _05271_ _05146_ _05253_ net1811 net1654 VPWR VGND sg13g2_a22oi_1
X_14103_ VPWR _00654_ net42 VGND sg13g2_inv_1
XFILLER_5_843 VPWR VGND sg13g2_decap_8
X_14034_ VPWR _00585_ net107 VGND sg13g2_inv_1
X_12295_ _06141_ _06139_ _06140_ VPWR VGND sg13g2_nand2_1
XFILLER_106_281 VPWR VGND sg13g2_decap_4
X_11246_ _05139_ _05144_ _05210_ VPWR VGND sg13g2_nor2_1
XFILLER_122_763 VPWR VGND sg13g2_decap_8
XFILLER_95_625 VPWR VGND sg13g2_fill_1
XFILLER_95_614 VPWR VGND sg13g2_decap_8
X_11177_ net1663 _05145_ _05146_ VPWR VGND sg13g2_nor2b_2
XFILLER_121_284 VPWR VGND sg13g2_fill_2
XFILLER_121_273 VPWR VGND sg13g2_decap_8
XFILLER_0_570 VPWR VGND sg13g2_decap_8
X_10128_ _04145_ _04138_ _04131_ _04210_ VPWR VGND sg13g2_nor3_2
XFILLER_110_969 VPWR VGND sg13g2_decap_8
XFILLER_94_157 VPWR VGND sg13g2_decap_8
X_14936_ _00737_ VGND VPWR _01456_ acc_sub.exp_mant_logic0.a\[4\] clknet_leaf_56_clk
+ sg13g2_dfrbpq_2
XFILLER_48_530 VPWR VGND sg13g2_decap_8
X_10059_ _04105_ VPWR _04147_ VGND _04144_ _04146_ sg13g2_o21ai_1
XFILLER_94_179 VPWR VGND sg13g2_fill_2
XFILLER_75_360 VPWR VGND sg13g2_decap_8
XFILLER_48_585 VPWR VGND sg13g2_decap_8
XFILLER_36_736 VPWR VGND sg13g2_decap_8
X_14867_ _00668_ VGND VPWR _01391_ fp16_sum_pipe.seg_reg0.q\[29\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_1
XFILLER_90_374 VPWR VGND sg13g2_fill_2
X_13818_ VPWR _00369_ net79 VGND sg13g2_inv_1
X_14798_ _00599_ VGND VPWR _01322_ acc_sum.exp_mant_logic0.a\[11\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_63_588 VPWR VGND sg13g2_fill_1
XFILLER_17_961 VPWR VGND sg13g2_decap_8
X_13749_ VPWR _00300_ net123 VGND sg13g2_inv_1
XFILLER_50_249 VPWR VGND sg13g2_decap_8
X_07270_ net1744 _01614_ _01638_ _01639_ VPWR VGND sg13g2_nand3_1
XFILLER_32_964 VPWR VGND sg13g2_decap_8
XFILLER_117_524 VPWR VGND sg13g2_decap_8
XFILLER_117_513 VPWR VGND sg13g2_fill_1
XFILLER_8_670 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_7_clk clknet_5_4__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
X_09911_ VPWR _04008_ _04007_ VGND sg13g2_inv_1
XFILLER_113_774 VPWR VGND sg13g2_decap_8
X_09842_ _03808_ _03804_ _03953_ VPWR VGND sg13g2_and2_1
XFILLER_99_986 VPWR VGND sg13g2_decap_8
X_09773_ _03889_ net1768 acc_sum.y\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_100_413 VPWR VGND sg13g2_decap_8
XFILLER_58_338 VPWR VGND sg13g2_decap_8
XFILLER_101_969 VPWR VGND sg13g2_decap_8
X_08724_ _02929_ VPWR _01329_ VGND net1815 _02928_ sg13g2_o21ai_1
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_96_1013 VPWR VGND sg13g2_fill_1
XFILLER_67_894 VPWR VGND sg13g2_fill_2
XFILLER_39_574 VPWR VGND sg13g2_decap_8
XFILLER_39_563 VPWR VGND sg13g2_decap_8
X_08655_ net1818 acc_sum.add_renorm0.mantisa\[8\] _02875_ VPWR VGND sg13g2_nor2_1
XFILLER_82_842 VPWR VGND sg13g2_fill_2
XFILLER_57_1008 VPWR VGND sg13g2_decap_4
XFILLER_26_246 VPWR VGND sg13g2_decap_8
X_07606_ _01914_ _01919_ _01920_ VPWR VGND sg13g2_nor2_1
X_08586_ _02809_ acc_sum.op_sign_logic0.mantisa_a\[9\] acc_sum.op_sign_logic0.mantisa_b\[9\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_82_886 VPWR VGND sg13g2_decap_4
XFILLER_26_257 VPWR VGND sg13g2_fill_2
XFILLER_26_268 VPWR VGND sg13g2_fill_2
X_07537_ _01856_ acc_sub.exp_mant_logic0.a\[10\] _01847_ _01779_ acc_sub.seg_reg0.q\[25\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_81_385 VPWR VGND sg13g2_fill_2
XFILLER_53_49 VPWR VGND sg13g2_fill_2
XFILLER_41_216 VPWR VGND sg13g2_decap_8
XFILLER_34_290 VPWR VGND sg13g2_decap_4
XFILLER_22_452 VPWR VGND sg13g2_decap_4
XFILLER_23_975 VPWR VGND sg13g2_decap_8
X_07468_ _01788_ _01790_ _01791_ VPWR VGND sg13g2_nor2_1
XFILLER_10_603 VPWR VGND sg13g2_decap_8
XFILLER_108_502 VPWR VGND sg13g2_decap_8
X_07399_ VPWR _01741_ acc_sub.exp_mant_logic0.a\[6\] VGND sg13g2_inv_1
X_09138_ net1787 _03227_ _03317_ VPWR VGND sg13g2_nor2_1
XFILLER_118_42 VPWR VGND sg13g2_decap_8
X_09069_ net1785 _03250_ _03253_ _03254_ VPWR VGND sg13g2_nor3_1
X_11100_ _02957_ _02959_ _02951_ _05071_ VPWR VGND _02963_ sg13g2_nand4_1
X_12080_ _05899_ _05925_ _05926_ VPWR VGND sg13g2_xor2_1
XFILLER_2_835 VPWR VGND sg13g2_decap_8
XFILLER_89_474 VPWR VGND sg13g2_decap_4
X_11031_ _05010_ _05009_ VPWR VGND _05007_ sg13g2_nand2b_2
XFILLER_1_345 VPWR VGND sg13g2_decap_8
XFILLER_104_785 VPWR VGND sg13g2_decap_8
XFILLER_76_135 VPWR VGND sg13g2_fill_1
XFILLER_92_628 VPWR VGND sg13g2_decap_8
X_12982_ _06750_ fpmul.seg_reg0.q\[15\] VPWR VGND sg13g2_inv_2
XFILLER_18_714 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_fill_2
XFILLER_57_382 VPWR VGND sg13g2_decap_8
XFILLER_45_522 VPWR VGND sg13g2_fill_1
X_11933_ VPWR _05799_ fpmul.seg_reg0.q\[35\] VGND sg13g2_inv_1
X_14721_ _00522_ VGND VPWR _01249_ fp16_res_pipe.exp_mant_logic0.a\[8\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
XFILLER_18_758 VPWR VGND sg13g2_fill_2
XFILLER_73_897 VPWR VGND sg13g2_decap_4
XFILLER_72_352 VPWR VGND sg13g2_decap_8
X_11864_ _05761_ _05573_ add_result\[7\] VPWR VGND sg13g2_nand2_1
X_14652_ _00453_ VGND VPWR _01180_ fp16_res_pipe.exp_mant_logic0.b\[5\] clknet_leaf_139_clk
+ sg13g2_dfrbpq_2
X_13603_ VPWR _00154_ net121 VGND sg13g2_inv_1
X_10815_ _04796_ _04802_ _04827_ VPWR VGND sg13g2_nor2_1
X_14583_ _00384_ VGND VPWR _01115_ fp16_sum_pipe.exp_mant_logic0.b\[10\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
X_11795_ _05697_ _05608_ _05622_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_430 VPWR VGND sg13g2_fill_1
XFILLER_32_249 VPWR VGND sg13g2_fill_1
X_13534_ VPWR _00085_ net85 VGND sg13g2_inv_1
XFILLER_9_412 VPWR VGND sg13g2_decap_4
XFILLER_13_463 VPWR VGND sg13g2_decap_8
XFILLER_14_986 VPWR VGND sg13g2_decap_8
X_10746_ _04759_ _04754_ _04758_ VPWR VGND sg13g2_nand2_2
X_13465_ _07112_ net1753 sipo.shift_reg\[1\] VPWR VGND sg13g2_nand2_1
X_10677_ _04690_ _04638_ _04615_ VPWR VGND sg13g2_nand2_1
XFILLER_127_855 VPWR VGND sg13g2_decap_8
XFILLER_126_343 VPWR VGND sg13g2_fill_1
X_13396_ _07074_ VPWR _00803_ VGND _05382_ net1696 sg13g2_o21ai_1
X_12347_ _06165_ _06192_ _06193_ VPWR VGND sg13g2_nor2_1
X_12278_ _06122_ _06123_ _06117_ _06124_ VPWR VGND sg13g2_nand3_1
XFILLER_4_161 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
X_11229_ _05194_ _05192_ VPWR VGND sg13g2_inv_2
X_14017_ VPWR _00568_ net22 VGND sg13g2_inv_1
XFILLER_122_571 VPWR VGND sg13g2_decap_8
XFILLER_96_934 VPWR VGND sg13g2_decap_8
XFILLER_67_124 VPWR VGND sg13g2_fill_1
XFILLER_4_98 VPWR VGND sg13g2_decap_8
XFILLER_110_766 VPWR VGND sg13g2_decap_8
XFILLER_67_135 VPWR VGND sg13g2_decap_8
XFILLER_67_168 VPWR VGND sg13g2_fill_1
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_48_360 VPWR VGND sg13g2_fill_2
X_14919_ _00720_ VGND VPWR _01439_ acc_sub.seg_reg0.q\[29\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_82_127 VPWR VGND sg13g2_fill_1
XFILLER_36_544 VPWR VGND sg13g2_decap_4
X_08440_ _02673_ VPWR _02674_ VGND fpdiv.divider0.divisor_reg\[8\] _02657_ sg13g2_o21ai_1
XFILLER_63_363 VPWR VGND sg13g2_decap_8
XFILLER_36_566 VPWR VGND sg13g2_decap_8
XFILLER_90_171 VPWR VGND sg13g2_decap_8
XFILLER_51_547 VPWR VGND sg13g2_fill_2
XFILLER_36_599 VPWR VGND sg13g2_decap_8
XFILLER_90_0 VPWR VGND sg13g2_decap_4
X_08371_ _02600_ _02613_ _02599_ _02614_ VPWR VGND sg13g2_nand3_1
XFILLER_17_1003 VPWR VGND sg13g2_decap_8
XFILLER_32_750 VPWR VGND sg13g2_fill_2
X_07322_ _01684_ VPWR _01685_ VGND _01561_ _01553_ sg13g2_o21ai_1
XFILLER_104_1006 VPWR VGND sg13g2_decap_8
XFILLER_20_934 VPWR VGND sg13g2_decap_8
X_07253_ VPWR _01623_ _01549_ VGND sg13g2_inv_1
X_07184_ VPWR _01556_ acc_sub.op_sign_logic0.mantisa_a\[3\] VGND sg13g2_inv_1
XFILLER_117_310 VPWR VGND sg13g2_fill_1
XFILLER_9_990 VPWR VGND sg13g2_decap_8
XFILLER_118_866 VPWR VGND sg13g2_decap_8
XFILLER_105_527 VPWR VGND sg13g2_decap_8
XFILLER_105_538 VPWR VGND sg13g2_fill_2
XFILLER_87_923 VPWR VGND sg13g2_decap_8
XFILLER_113_582 VPWR VGND sg13g2_fill_1
X_09825_ VGND VPWR _03851_ _03628_ _03937_ _03858_ sg13g2_a21oi_1
XFILLER_101_711 VPWR VGND sg13g2_fill_2
XFILLER_86_400 VPWR VGND sg13g2_decap_4
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_58_135 VPWR VGND sg13g2_decap_8
X_09756_ VPWR _03872_ _03871_ VGND sg13g2_inv_1
XFILLER_100_265 VPWR VGND sg13g2_fill_2
XFILLER_73_116 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_fill_1
XFILLER_104_55 VPWR VGND sg13g2_fill_1
XFILLER_100_287 VPWR VGND sg13g2_decap_8
X_09687_ _03802_ VPWR _03803_ VGND acc_sum.add_renorm0.mantisa\[11\] _02928_ sg13g2_o21ai_1
X_08707_ _02803_ _02841_ _02842_ _02919_ VPWR VGND sg13g2_nor3_1
XFILLER_54_330 VPWR VGND sg13g2_fill_2
XFILLER_27_522 VPWR VGND sg13g2_decap_4
X_08638_ _02860_ _02840_ _02859_ VPWR VGND sg13g2_xnor2_1
XFILLER_54_352 VPWR VGND sg13g2_decap_8
XFILLER_15_706 VPWR VGND sg13g2_fill_2
XFILLER_120_21 VPWR VGND sg13g2_decap_8
XFILLER_70_834 VPWR VGND sg13g2_fill_2
XFILLER_14_238 VPWR VGND sg13g2_decap_4
X_08569_ VPWR VGND _02792_ _02730_ _02787_ _02732_ _02793_ _02733_ sg13g2_a221oi_1
Xfanout20 net24 net20 VPWR VGND sg13g2_buf_2
Xfanout31 net39 net31 VPWR VGND sg13g2_buf_2
XFILLER_120_98 VPWR VGND sg13g2_decap_8
XFILLER_80_25 VPWR VGND sg13g2_fill_1
Xfanout64 net67 net64 VPWR VGND sg13g2_buf_1
Xfanout53 net55 net53 VPWR VGND sg13g2_buf_1
Xfanout42 net47 net42 VPWR VGND sg13g2_buf_2
X_10600_ VPWR _04613_ fp16_res_pipe.add_renorm0.mantisa\[6\] VGND sg13g2_inv_1
X_11580_ VPWR _05485_ _05484_ VGND sg13g2_inv_1
XFILLER_22_260 VPWR VGND sg13g2_decap_8
XFILLER_23_783 VPWR VGND sg13g2_fill_1
XFILLER_109_800 VPWR VGND sg13g2_decap_8
Xfanout97 net100 net97 VPWR VGND sg13g2_buf_2
Xfanout75 net76 net75 VPWR VGND sg13g2_buf_2
Xfanout86 net93 net86 VPWR VGND sg13g2_buf_2
XFILLER_7_916 VPWR VGND sg13g2_decap_8
X_10531_ _04571_ _04569_ _04570_ _04477_ net1737 VPWR VGND sg13g2_a22oi_1
XFILLER_11_945 VPWR VGND sg13g2_decap_8
X_13250_ _06974_ net1743 sipo.word\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_13_63 VPWR VGND sg13g2_decap_8
XFILLER_89_23 VPWR VGND sg13g2_fill_2
X_12201_ VPWR _06047_ _06045_ VGND sg13g2_inv_1
X_10462_ VPWR _04510_ _04509_ VGND sg13g2_inv_1
XFILLER_10_488 VPWR VGND sg13g2_decap_4
XFILLER_89_45 VPWR VGND sg13g2_decap_8
X_13181_ _06922_ net1715 sipo.word\[10\] VPWR VGND sg13g2_nand2_1
X_10393_ VPWR _04443_ _04442_ VGND sg13g2_inv_1
XFILLER_124_858 VPWR VGND sg13g2_decap_8
XFILLER_123_346 VPWR VGND sg13g2_decap_8
XFILLER_89_89 VPWR VGND sg13g2_decap_8
X_12132_ VPWR _05978_ _05977_ VGND sg13g2_inv_1
XFILLER_2_632 VPWR VGND sg13g2_decap_8
XFILLER_123_379 VPWR VGND sg13g2_fill_2
XFILLER_96_219 VPWR VGND sg13g2_fill_1
X_12063_ VPWR _05909_ _05883_ VGND sg13g2_inv_1
XFILLER_78_956 VPWR VGND sg13g2_fill_2
XFILLER_78_923 VPWR VGND sg13g2_decap_4
X_11014_ acc_sum.reg1en.q\[0\] _04993_ VPWR VGND sg13g2_inv_4
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_78_967 VPWR VGND sg13g2_fill_2
XFILLER_93_926 VPWR VGND sg13g2_decap_8
XFILLER_65_628 VPWR VGND sg13g2_decap_4
XFILLER_49_168 VPWR VGND sg13g2_fill_1
XFILLER_37_308 VPWR VGND sg13g2_decap_4
X_12965_ _06736_ net1717 _00006_ VPWR VGND sg13g2_nand2_1
X_14704_ _00505_ VGND VPWR _01232_ acc_sum.y\[7\] clknet_leaf_23_clk sg13g2_dfrbpq_1
X_11916_ _05788_ net1882 fpmul.reg_a_out\[2\] VPWR VGND sg13g2_nand2_1
X_12896_ VGND VPWR net1936 add_result\[6\] _06672_ net1950 sg13g2_a21oi_1
XFILLER_61_878 VPWR VGND sg13g2_decap_4
XFILLER_54_81 VPWR VGND sg13g2_decap_4
X_14635_ _00436_ VGND VPWR _01167_ fp16_sum_pipe.add_renorm0.mantisa\[6\] clknet_leaf_108_clk
+ sg13g2_dfrbpq_2
X_11847_ _05648_ _05744_ _05745_ VPWR VGND _05743_ sg13g2_nand3b_1
X_14566_ _00367_ VGND VPWR _01102_ acc_sum.seg_reg0.q\[29\] clknet_leaf_25_clk sg13g2_dfrbpq_1
X_11778_ _05681_ _05644_ _05628_ VPWR VGND sg13g2_nand2_1
XFILLER_20_219 VPWR VGND sg13g2_decap_8
XFILLER_119_608 VPWR VGND sg13g2_fill_1
X_13517_ VPWR _00068_ net84 VGND sg13g2_inv_1
X_10729_ _04670_ _04726_ _04742_ VPWR VGND sg13g2_nor2_2
X_14497_ _00298_ VGND VPWR _01033_ fpdiv.divider0.divisor\[8\] clknet_leaf_85_clk
+ sg13g2_dfrbpq_1
XFILLER_9_275 VPWR VGND sg13g2_decap_8
XFILLER_9_286 VPWR VGND sg13g2_fill_2
XFILLER_86_1001 VPWR VGND sg13g2_decap_8
Xclkload12 clknet_5_25__leaf_clk clkload12/X VPWR VGND sg13g2_buf_8
Xclkload34 clknet_leaf_4_clk clkload34/Y VPWR VGND sg13g2_inv_4
X_13448_ _07103_ VPWR _00780_ VGND _06920_ net1754 sg13g2_o21ai_1
Xclkload23 clkload23/Y clknet_leaf_136_clk VPWR VGND sg13g2_inv_8
XFILLER_126_140 VPWR VGND sg13g2_decap_8
XFILLER_86_1012 VPWR VGND sg13g2_fill_2
Xclkload78 clkload78/Y clknet_leaf_55_clk VPWR VGND sg13g2_inv_8
Xclkload67 clknet_leaf_26_clk clkload67/Y VPWR VGND sg13g2_inv_4
X_13379_ _07066_ _07055_ sipo.word\[9\] VPWR VGND sg13g2_nand2_1
Xclkload56 clkload56/Y clknet_leaf_124_clk VPWR VGND sg13g2_inv_2
Xclkload45 clkload45/Y clknet_leaf_118_clk VPWR VGND sg13g2_inv_8
XFILLER_115_858 VPWR VGND sg13g2_decap_8
Xclkload89 clknet_leaf_44_clk clkload89/Y VPWR VGND sg13g2_inv_4
XFILLER_5_492 VPWR VGND sg13g2_decap_8
XFILLER_88_709 VPWR VGND sg13g2_decap_8
XFILLER_69_912 VPWR VGND sg13g2_fill_1
XFILLER_69_901 VPWR VGND sg13g2_fill_1
X_07940_ VPWR _02215_ _02214_ VGND sg13g2_inv_1
XFILLER_95_230 VPWR VGND sg13g2_fill_1
X_07871_ _02162_ VPWR _01408_ VGND net1887 _01789_ sg13g2_o21ai_1
XFILLER_69_956 VPWR VGND sg13g2_decap_8
X_09610_ _03692_ _03697_ _03727_ VPWR VGND sg13g2_nor2_1
XFILLER_28_308 VPWR VGND sg13g2_fill_2
X_09541_ _03628_ _03640_ _03644_ _03658_ VPWR VGND sg13g2_nand3_1
XFILLER_84_959 VPWR VGND sg13g2_decap_8
XFILLER_92_981 VPWR VGND sg13g2_decap_8
XFILLER_52_812 VPWR VGND sg13g2_fill_1
XFILLER_37_875 VPWR VGND sg13g2_decap_8
XFILLER_36_396 VPWR VGND sg13g2_fill_1
XFILLER_36_374 VPWR VGND sg13g2_decap_8
X_09472_ VPWR _03599_ fp16_res_pipe.exp_mant_logic0.a\[9\] VGND sg13g2_inv_1
X_08423_ VPWR _02657_ fpdiv.divider0.remainder_reg\[8\] VGND sg13g2_inv_1
XFILLER_12_709 VPWR VGND sg13g2_decap_8
X_08354_ instr\[15\] instr\[14\] instr\[13\] instr\[12\] _02597_ VPWR VGND sg13g2_nor4_1
XFILLER_11_219 VPWR VGND sg13g2_decap_8
X_07305_ _01668_ _01670_ _01667_ _01482_ VPWR VGND sg13g2_nand3_1
Xclkload6 clknet_5_13__leaf_clk clkload6/X VPWR VGND sg13g2_buf_8
XFILLER_50_28 VPWR VGND sg13g2_decap_8
X_08285_ _02530_ _02532_ _02533_ VPWR VGND sg13g2_nor2_1
X_07236_ _01606_ VPWR _01607_ VGND _01531_ _01533_ sg13g2_o21ai_1
XFILLER_118_652 VPWR VGND sg13g2_decap_8
XFILLER_30_1011 VPWR VGND sg13g2_fill_2
X_07167_ VPWR _01539_ acc_sub.op_sign_logic0.mantisa_b\[4\] VGND sg13g2_inv_1
XFILLER_117_140 VPWR VGND sg13g2_decap_8
XFILLER_78_208 VPWR VGND sg13g2_fill_2
XFILLER_120_327 VPWR VGND sg13g2_fill_1
XFILLER_120_305 VPWR VGND sg13g2_fill_2
XFILLER_115_21 VPWR VGND sg13g2_decap_8
XFILLER_99_591 VPWR VGND sg13g2_fill_1
XFILLER_99_580 VPWR VGND sg13g2_decap_8
XFILLER_59_411 VPWR VGND sg13g2_fill_1
XFILLER_113_390 VPWR VGND sg13g2_decap_4
X_09808_ _03921_ _03836_ _03871_ VPWR VGND sg13g2_xnor2_1
XFILLER_87_775 VPWR VGND sg13g2_fill_1
XFILLER_75_948 VPWR VGND sg13g2_decap_8
XFILLER_59_477 VPWR VGND sg13g2_decap_8
XFILLER_47_639 VPWR VGND sg13g2_decap_8
XFILLER_47_606 VPWR VGND sg13g2_fill_2
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_115_98 VPWR VGND sg13g2_decap_8
X_09739_ _03853_ _03854_ _03855_ VPWR VGND sg13g2_and2_1
XFILLER_86_296 VPWR VGND sg13g2_fill_2
XFILLER_28_831 VPWR VGND sg13g2_fill_1
XFILLER_27_341 VPWR VGND sg13g2_fill_1
XFILLER_83_981 VPWR VGND sg13g2_decap_8
X_12750_ fpmul.reg_b_out\[7\] fp16_res_pipe.x2\[7\] net1955 _00917_ VPWR VGND sg13g2_mux2_1
XFILLER_91_46 VPWR VGND sg13g2_decap_4
X_12681_ _06493_ _06462_ _06418_ VPWR VGND sg13g2_nand2_1
XFILLER_43_867 VPWR VGND sg13g2_decap_8
XFILLER_15_558 VPWR VGND sg13g2_decap_8
X_14420_ _00221_ VGND VPWR _00959_ fpmul.seg_reg0.q\[5\] clknet_leaf_78_clk sg13g2_dfrbpq_1
X_11632_ VPWR _05537_ _05536_ VGND sg13g2_inv_1
XFILLER_30_517 VPWR VGND sg13g2_fill_1
XFILLER_30_528 VPWR VGND sg13g2_decap_8
X_14351_ _00152_ VGND VPWR _00893_ fpmul.reg_p_out\[15\] clknet_leaf_90_clk sg13g2_dfrbpq_1
XFILLER_24_84 VPWR VGND sg13g2_decap_8
XFILLER_30_539 VPWR VGND sg13g2_fill_1
X_13302_ _07014_ sipo.word\[2\] VPWR VGND sg13g2_inv_2
X_11563_ _05468_ _05457_ _05459_ VPWR VGND sg13g2_nand2_1
X_14282_ _00083_ VGND VPWR _00833_ fp16_res_pipe.x2\[15\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_10514_ VGND VPWR _04555_ net1848 _01166_ _04556_ sg13g2_a21oi_1
XFILLER_7_746 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_fill_1
XFILLER_10_274 VPWR VGND sg13g2_decap_4
X_11494_ _05399_ net1840 fp16_sum_pipe.add_renorm0.mantisa\[8\] VPWR VGND sg13g2_nand2_1
X_13233_ _02611_ _02607_ _02600_ _06958_ VPWR VGND sg13g2_nand3_1
XFILLER_6_267 VPWR VGND sg13g2_decap_8
X_10445_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[8\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[8\]
+ net1736 _04494_ VPWR VGND sg13g2_nand3_1
XFILLER_108_173 VPWR VGND sg13g2_decap_4
X_13164_ _06910_ net1713 sipo.word\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_123_154 VPWR VGND sg13g2_decap_8
XFILLER_112_817 VPWR VGND sg13g2_decap_8
XFILLER_97_506 VPWR VGND sg13g2_fill_2
X_12115_ _05961_ _05958_ _05960_ VPWR VGND sg13g2_xnor2_1
X_10376_ _04426_ _04424_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_3_952 VPWR VGND sg13g2_decap_8
X_13095_ _06855_ VPWR _00885_ VGND net1862 _06666_ sg13g2_o21ai_1
XFILLER_2_451 VPWR VGND sg13g2_decap_8
XFILLER_77_241 VPWR VGND sg13g2_fill_1
X_12046_ _05892_ _05890_ _05891_ VPWR VGND sg13g2_nand2_1
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_120_883 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_93_745 VPWR VGND sg13g2_fill_1
XFILLER_77_296 VPWR VGND sg13g2_decap_8
XFILLER_37_138 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
X_13997_ VPWR _00548_ net10 VGND sg13g2_inv_1
X_12948_ _06720_ _06716_ _06719_ _06533_ net1948 VPWR VGND sg13g2_a22oi_1
XFILLER_46_694 VPWR VGND sg13g2_decap_8
XFILLER_34_845 VPWR VGND sg13g2_decap_8
X_12879_ _06656_ VPWR _06657_ VGND fpmul.reg1en.d\[0\] _06654_ sg13g2_o21ai_1
XFILLER_61_653 VPWR VGND sg13g2_fill_1
XFILLER_45_182 VPWR VGND sg13g2_decap_8
XFILLER_34_856 VPWR VGND sg13g2_fill_2
X_14618_ _00419_ VGND VPWR _01150_ fp16_sum_pipe.exp_mant_logic0.a\[13\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_1
XFILLER_21_528 VPWR VGND sg13g2_decap_8
XFILLER_60_196 VPWR VGND sg13g2_decap_8
XFILLER_21_539 VPWR VGND sg13g2_fill_2
XFILLER_119_405 VPWR VGND sg13g2_decap_4
X_14549_ _00350_ VGND VPWR _01085_ acc_sum.op_sign_logic0.mantisa_a\[1\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
Xclkload112 VPWR clkload112/Y clknet_leaf_67_clk VGND sg13g2_inv_1
Xclkload101 clkload101/Y clknet_leaf_75_clk VPWR VGND sg13g2_inv_2
X_08070_ _02336_ _02220_ _02214_ VPWR VGND sg13g2_nand2_1
XFILLER_115_600 VPWR VGND sg13g2_decap_8
Xplace1902 net1900 net1902 VPWR VGND sg13g2_buf_1
XFILLER_115_644 VPWR VGND sg13g2_decap_8
Xplace1946 net1944 net1946 VPWR VGND sg13g2_buf_2
Xplace1935 net1923 net1935 VPWR VGND sg13g2_buf_2
XFILLER_53_0 VPWR VGND sg13g2_decap_8
Xplace1924 net1923 net1924 VPWR VGND sg13g2_buf_2
Xplace1913 net1912 net1913 VPWR VGND sg13g2_buf_2
XFILLER_6_790 VPWR VGND sg13g2_decap_4
XFILLER_114_154 VPWR VGND sg13g2_decap_8
Xplace1957 net1954 net1957 VPWR VGND sg13g2_buf_2
X_08972_ _03158_ _03085_ _03084_ VPWR VGND sg13g2_nand2_1
X_07923_ fp16_sum_pipe.exp_mant_logic0.b\[12\] _02197_ _02198_ VPWR VGND sg13g2_nor2_1
X_07854_ _02149_ net1779 acc_sub.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_57_926 VPWR VGND sg13g2_decap_8
XFILLER_111_894 VPWR VGND sg13g2_decap_8
XFILLER_83_211 VPWR VGND sg13g2_decap_8
XFILLER_68_296 VPWR VGND sg13g2_decap_4
XFILLER_57_959 VPWR VGND sg13g2_decap_8
XFILLER_28_116 VPWR VGND sg13g2_fill_2
X_07785_ _02085_ _02084_ net1640 VPWR VGND sg13g2_nand2_1
XFILLER_45_28 VPWR VGND sg13g2_decap_8
X_09524_ VPWR _03641_ _03640_ VGND sg13g2_inv_1
XFILLER_65_981 VPWR VGND sg13g2_decap_8
XFILLER_43_119 VPWR VGND sg13g2_decap_8
XFILLER_52_653 VPWR VGND sg13g2_fill_1
XFILLER_52_642 VPWR VGND sg13g2_fill_1
X_09455_ fp16_res_pipe.exp_mant_logic0.a\[15\] net1911 _03588_ VPWR VGND sg13g2_nor2_1
XFILLER_101_56 VPWR VGND sg13g2_decap_8
XFILLER_80_984 VPWR VGND sg13g2_decap_8
X_08406_ _02642_ _02589_ state\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_52_664 VPWR VGND sg13g2_decap_8
XFILLER_51_141 VPWR VGND sg13g2_fill_2
XFILLER_12_528 VPWR VGND sg13g2_decap_8
XFILLER_25_889 VPWR VGND sg13g2_decap_8
XFILLER_51_196 VPWR VGND sg13g2_decap_8
X_09386_ net1738 _03471_ _03533_ _03534_ VPWR VGND sg13g2_nand3_1
X_08337_ _02582_ sipo.word_ready VPWR VGND sg13g2_inv_2
X_08268_ _02517_ net1657 fp16_sum_pipe.exp_mant_logic0.b\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_20_594 VPWR VGND sg13g2_decap_8
XFILLER_119_961 VPWR VGND sg13g2_decap_8
X_07219_ _01500_ _01590_ _01591_ VPWR VGND sg13g2_nor2b_2
X_08199_ _02456_ net1774 fp16_sum_pipe.op_sign_logic0.mantisa_a\[0\] VPWR VGND sg13g2_nand2_1
X_10230_ _04302_ _04175_ _04303_ VPWR VGND sg13g2_nor2_1
XFILLER_106_677 VPWR VGND sg13g2_decap_8
XFILLER_10_42 VPWR VGND sg13g2_decap_8
XFILLER_126_42 VPWR VGND sg13g2_decap_8
XFILLER_117_1005 VPWR VGND sg13g2_decap_8
XFILLER_105_176 VPWR VGND sg13g2_decap_8
X_10161_ _04242_ net1764 fp16_res_pipe.op_sign_logic0.mantisa_a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_59_230 VPWR VGND sg13g2_decap_8
XFILLER_0_933 VPWR VGND sg13g2_decap_8
X_10092_ _04175_ _04177_ VPWR VGND sg13g2_inv_4
XFILLER_120_168 VPWR VGND sg13g2_decap_8
XFILLER_86_79 VPWR VGND sg13g2_decap_4
X_13920_ VPWR _00471_ net5 VGND sg13g2_inv_1
XFILLER_101_393 VPWR VGND sg13g2_decap_8
XFILLER_19_127 VPWR VGND sg13g2_decap_8
XFILLER_75_778 VPWR VGND sg13g2_fill_2
X_13851_ VPWR _00402_ net30 VGND sg13g2_inv_1
X_13782_ VPWR _00333_ net126 VGND sg13g2_inv_1
X_12802_ VPWR _06586_ fpmul.reg_p_out\[14\] VGND sg13g2_inv_1
X_10994_ _04983_ fp16_res_pipe.x2\[7\] net1933 VPWR VGND sg13g2_nand2_1
XFILLER_34_119 VPWR VGND sg13g2_decap_8
XFILLER_16_834 VPWR VGND sg13g2_fill_2
X_12733_ VPWR _06536_ div_result\[1\] VGND sg13g2_inv_1
XFILLER_16_889 VPWR VGND sg13g2_decap_8
X_12664_ _06479_ VPWR _06480_ VGND net1735 _06477_ sg13g2_o21ai_1
XFILLER_70_494 VPWR VGND sg13g2_decap_4
X_14403_ _00204_ VGND VPWR _00942_ fpmul.reg_a_out\[0\] clknet_leaf_103_clk sg13g2_dfrbpq_1
XFILLER_43_697 VPWR VGND sg13g2_decap_8
XFILLER_42_196 VPWR VGND sg13g2_fill_2
XFILLER_15_388 VPWR VGND sg13g2_fill_1
XFILLER_89_9 VPWR VGND sg13g2_fill_1
X_12595_ _06410_ _06409_ _06411_ VPWR VGND sg13g2_xor2_1
X_11615_ fp16_sum_pipe.add_renorm0.mantisa\[1\] _05519_ _05412_ _05520_ VPWR VGND
+ sg13g2_nor3_1
X_14334_ _00135_ VGND VPWR _00876_ piso.tx_bit_counter\[3\] clknet_leaf_86_clk sg13g2_dfrbpq_1
X_11546_ VPWR _05451_ fp16_sum_pipe.add_renorm0.mantisa\[9\] VGND sg13g2_inv_1
XFILLER_116_419 VPWR VGND sg13g2_fill_1
X_14265_ _00066_ VGND VPWR _00816_ acc_sub.x2\[14\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_125_942 VPWR VGND sg13g2_decap_8
X_11477_ _05390_ VPWR _01037_ VGND net1937 _05389_ sg13g2_o21ai_1
X_13216_ _06944_ _06943_ _00853_ VPWR VGND sg13g2_nor2_1
X_14196_ VPWR _00747_ net91 VGND sg13g2_inv_1
X_10428_ _04477_ _04475_ _04476_ VPWR VGND sg13g2_nand2_1
XFILLER_124_485 VPWR VGND sg13g2_decap_8
XFILLER_112_625 VPWR VGND sg13g2_decap_8
XFILLER_98_826 VPWR VGND sg13g2_decap_8
XFILLER_97_314 VPWR VGND sg13g2_decap_8
X_13147_ _06895_ _06566_ net4 VPWR VGND sg13g2_nand2_1
X_10359_ VPWR _04409_ _04408_ VGND sg13g2_inv_1
XFILLER_124_496 VPWR VGND sg13g2_fill_1
X_13078_ _06844_ _06843_ _06815_ VPWR VGND sg13g2_nand2_1
XFILLER_66_712 VPWR VGND sg13g2_decap_8
X_12029_ _05876_ fpmul.reg1en.q\[0\] VPWR VGND sg13g2_inv_2
XFILLER_65_222 VPWR VGND sg13g2_fill_2
XFILLER_65_211 VPWR VGND sg13g2_fill_1
XFILLER_65_200 VPWR VGND sg13g2_fill_1
XFILLER_65_266 VPWR VGND sg13g2_decap_8
XFILLER_65_255 VPWR VGND sg13g2_fill_2
X_07570_ VPWR _01884_ _01883_ VGND sg13g2_inv_1
XFILLER_81_748 VPWR VGND sg13g2_fill_2
XFILLER_81_737 VPWR VGND sg13g2_decap_8
XFILLER_65_288 VPWR VGND sg13g2_fill_1
XFILLER_47_981 VPWR VGND sg13g2_fill_2
XFILLER_18_182 VPWR VGND sg13g2_decap_8
X_09240_ VPWR _03394_ fp16_res_pipe.op_sign_logic0.mantisa_a\[5\] VGND sg13g2_inv_1
XFILLER_21_325 VPWR VGND sg13g2_fill_2
XFILLER_22_848 VPWR VGND sg13g2_decap_8
X_09171_ VPWR _03337_ acc_sum.exp_mant_logic0.b\[10\] VGND sg13g2_inv_1
XFILLER_21_369 VPWR VGND sg13g2_decap_8
XFILLER_119_224 VPWR VGND sg13g2_decap_8
XFILLER_108_909 VPWR VGND sg13g2_decap_8
X_08122_ _02376_ _02381_ _02383_ _02384_ VPWR VGND sg13g2_nor3_1
XFILLER_30_892 VPWR VGND sg13g2_decap_8
X_08053_ VPWR _02319_ _02220_ VGND sg13g2_inv_1
Xplace1710 _04654_ net1710 VPWR VGND sg13g2_buf_2
XFILLER_116_975 VPWR VGND sg13g2_decap_8
Xplace1743 net1742 net1743 VPWR VGND sg13g2_buf_1
XFILLER_89_815 VPWR VGND sg13g2_decap_8
Xplace1732 _06559_ net1732 VPWR VGND sg13g2_buf_2
Xplace1721 _07076_ net1721 VPWR VGND sg13g2_buf_2
Xplace1754 net1751 net1754 VPWR VGND sg13g2_buf_2
Xplace1787 acc_sub.seg_reg1.q\[21\] net1787 VPWR VGND sg13g2_buf_2
Xplace1776 net1775 net1776 VPWR VGND sg13g2_buf_2
Xplace1765 _03988_ net1765 VPWR VGND sg13g2_buf_2
Xplace1798 net1797 net1798 VPWR VGND sg13g2_buf_1
X_08955_ _03141_ _03140_ acc_sub.add_renorm0.exp\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_103_647 VPWR VGND sg13g2_fill_1
XFILLER_102_124 VPWR VGND sg13g2_decap_4
XFILLER_102_113 VPWR VGND sg13g2_fill_2
XFILLER_102_179 VPWR VGND sg13g2_fill_1
XFILLER_5_1004 VPWR VGND sg13g2_decap_8
X_08886_ _03072_ _01490_ _03073_ VPWR VGND sg13g2_and2_1
XFILLER_111_691 VPWR VGND sg13g2_decap_4
XFILLER_99_1000 VPWR VGND sg13g2_decap_8
XFILLER_84_520 VPWR VGND sg13g2_fill_2
XFILLER_29_414 VPWR VGND sg13g2_fill_2
X_07837_ _02133_ _01959_ acc_sub.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_nand2_1
X_07768_ _02068_ _02069_ _02067_ _02070_ VPWR VGND sg13g2_nand3_1
XFILLER_72_737 VPWR VGND sg13g2_fill_1
XFILLER_44_428 VPWR VGND sg13g2_fill_1
XFILLER_16_108 VPWR VGND sg13g2_decap_8
XFILLER_112_77 VPWR VGND sg13g2_decap_8
X_09507_ _03620_ _03623_ _03624_ VPWR VGND sg13g2_nor2_1
XFILLER_71_258 VPWR VGND sg13g2_decap_8
XFILLER_53_962 VPWR VGND sg13g2_fill_2
XFILLER_53_951 VPWR VGND sg13g2_decap_4
XFILLER_72_48 VPWR VGND sg13g2_fill_1
XFILLER_40_612 VPWR VGND sg13g2_decap_8
XFILLER_13_815 VPWR VGND sg13g2_decap_4
XFILLER_24_141 VPWR VGND sg13g2_decap_4
XFILLER_52_483 VPWR VGND sg13g2_decap_8
X_09438_ _03577_ VPWR _01263_ VGND net1834 _03576_ sg13g2_o21ai_1
X_09369_ _03518_ VPWR _03519_ VGND _03516_ _03517_ sg13g2_o21ai_1
X_11400_ _05344_ VPWR _01068_ VGND _05342_ fpdiv.divider0.en_r sg13g2_o21ai_1
X_12380_ _06225_ VPWR _06226_ VGND _05891_ _06015_ sg13g2_o21ai_1
X_11331_ _05286_ net1634 _05285_ VPWR VGND sg13g2_nand2_1
XFILLER_125_238 VPWR VGND sg13g2_decap_8
XFILLER_21_63 VPWR VGND sg13g2_decap_8
XFILLER_107_964 VPWR VGND sg13g2_decap_8
X_11262_ _05221_ _05224_ _05225_ VPWR VGND sg13g2_nor2_1
X_14050_ VPWR _00601_ net22 VGND sg13g2_inv_1
X_11193_ _05122_ _05112_ net1663 _05161_ VPWR VGND sg13g2_nor3_2
X_13001_ _06769_ fpmul.seg_reg0.q\[15\] fpmul.seg_reg0.q\[13\] VPWR VGND sg13g2_nand2_1
X_10213_ _01198_ _04286_ _04287_ VPWR VGND sg13g2_nand2_1
XFILLER_122_945 VPWR VGND sg13g2_decap_8
X_10144_ _04225_ _04224_ net1746 VPWR VGND sg13g2_nand2_1
X_14952_ _00753_ VGND VPWR _01472_ acc_sub.add_renorm0.exp\[4\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_2
XFILLER_87_380 VPWR VGND sg13g2_decap_4
XFILLER_75_520 VPWR VGND sg13g2_decap_4
X_10075_ _04162_ net1637 _04161_ VPWR VGND sg13g2_nand2_1
XFILLER_101_190 VPWR VGND sg13g2_decap_4
X_14883_ _00684_ VGND VPWR _01403_ acc_sub.exp_mant_logic0.b\[9\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
X_13903_ VPWR _00454_ net7 VGND sg13g2_inv_1
XFILLER_90_501 VPWR VGND sg13g2_fill_1
XFILLER_75_597 VPWR VGND sg13g2_decap_8
XFILLER_62_203 VPWR VGND sg13g2_fill_2
X_13834_ VPWR _00385_ net14 VGND sg13g2_inv_1
XFILLER_90_545 VPWR VGND sg13g2_decap_4
XFILLER_90_534 VPWR VGND sg13g2_fill_1
XFILLER_62_247 VPWR VGND sg13g2_decap_8
XFILLER_16_642 VPWR VGND sg13g2_fill_1
X_13765_ VPWR _00316_ net129 VGND sg13g2_inv_1
X_10977_ _04975_ _04772_ fp16_res_pipe.y\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_94_7 VPWR VGND sg13g2_decap_8
X_12716_ _06522_ _06450_ _06437_ VPWR VGND sg13g2_nand2_1
XFILLER_70_280 VPWR VGND sg13g2_decap_8
X_13696_ VPWR _00247_ net61 VGND sg13g2_inv_1
XFILLER_43_483 VPWR VGND sg13g2_decap_8
XFILLER_15_196 VPWR VGND sg13g2_decap_8
X_12647_ _06418_ _06462_ _06463_ VPWR VGND sg13g2_nor2_1
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_30_188 VPWR VGND sg13g2_fill_1
X_12578_ _06392_ _06389_ _06393_ _06394_ VPWR VGND sg13g2_a21o_1
XFILLER_8_874 VPWR VGND sg13g2_decap_8
XFILLER_117_739 VPWR VGND sg13g2_decap_8
X_14317_ _00118_ VGND VPWR _00860_ sipo.word\[5\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_7_373 VPWR VGND sg13g2_fill_2
X_11529_ VGND VPWR _05433_ _05434_ _05432_ _05431_ sg13g2_a21oi_2
X_14248_ _00049_ VGND VPWR _00799_ instr\[13\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_7_98 VPWR VGND sg13g2_decap_8
X_14179_ VPWR _00730_ net127 VGND sg13g2_inv_1
XFILLER_113_956 VPWR VGND sg13g2_decap_8
XFILLER_112_444 VPWR VGND sg13g2_decap_8
XFILLER_86_807 VPWR VGND sg13g2_decap_8
XFILLER_39_701 VPWR VGND sg13g2_fill_1
X_08740_ _02940_ acc\[12\] net1901 VPWR VGND sg13g2_nand2_1
X_08671_ VGND VPWR _02887_ net1818 _01341_ _02888_ sg13g2_a21oi_1
XFILLER_66_542 VPWR VGND sg13g2_fill_2
XFILLER_38_244 VPWR VGND sg13g2_decap_8
XFILLER_16_0 VPWR VGND sg13g2_decap_8
XFILLER_27_918 VPWR VGND sg13g2_decap_8
X_07622_ _01880_ _01817_ _01936_ VPWR VGND sg13g2_nor2_1
XFILLER_54_726 VPWR VGND sg13g2_fill_2
XFILLER_39_789 VPWR VGND sg13g2_decap_8
XFILLER_53_247 VPWR VGND sg13g2_decap_8
XFILLER_53_225 VPWR VGND sg13g2_decap_4
X_07553_ _01864_ _01865_ _01866_ _01868_ VGND VPWR _01867_ sg13g2_nor4_2
X_07484_ acc_sub.exp_mant_logic0.b\[9\] _01735_ _01807_ VPWR VGND sg13g2_nor2_1
XFILLER_35_995 VPWR VGND sg13g2_decap_8
XFILLER_10_807 VPWR VGND sg13g2_decap_8
X_09223_ VPWR _03377_ _03376_ VGND sg13g2_inv_1
XFILLER_21_133 VPWR VGND sg13g2_fill_2
X_09154_ _03326_ net1773 acc_sub.y\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_50_998 VPWR VGND sg13g2_decap_8
XFILLER_108_717 VPWR VGND sg13g2_fill_2
X_08105_ _02369_ fp16_sum_pipe.exp_mant_logic0.a\[4\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[7\]
+ net1776 VPWR VGND sg13g2_a22oi_1
X_09085_ net1785 _03266_ _03268_ _03269_ VPWR VGND sg13g2_nor3_1
XFILLER_107_216 VPWR VGND sg13g2_fill_1
XFILLER_107_205 VPWR VGND sg13g2_decap_8
X_08036_ VGND VPWR _02289_ _02245_ _02302_ _02301_ sg13g2_a21oi_1
XFILLER_116_772 VPWR VGND sg13g2_decap_8
XFILLER_104_901 VPWR VGND sg13g2_decap_8
XFILLER_107_55 VPWR VGND sg13g2_decap_8
XFILLER_103_422 VPWR VGND sg13g2_decap_8
XFILLER_1_527 VPWR VGND sg13g2_decap_8
XFILLER_104_978 VPWR VGND sg13g2_decap_8
X_09987_ _04075_ VPWR _01212_ VGND net1831 _03444_ sg13g2_o21ai_1
X_08938_ VGND VPWR _03124_ _03125_ net1787 _03122_ sg13g2_a21oi_2
XFILLER_103_499 VPWR VGND sg13g2_fill_1
XFILLER_88_199 VPWR VGND sg13g2_fill_1
X_08869_ _03056_ _03024_ _01707_ acc_sub.add_renorm0.mantisa\[3\] _02985_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_123_21 VPWR VGND sg13g2_decap_8
XFILLER_83_25 VPWR VGND sg13g2_decap_4
X_10900_ net1772 _04907_ _04909_ _04910_ VPWR VGND sg13g2_nor3_1
XFILLER_123_98 VPWR VGND sg13g2_decap_8
X_11880_ _02645_ _05768_ _05769_ VPWR VGND sg13g2_nor2_1
XFILLER_17_439 VPWR VGND sg13g2_decap_8
XFILLER_26_940 VPWR VGND sg13g2_decap_8
XFILLER_72_578 VPWR VGND sg13g2_decap_8
XFILLER_44_258 VPWR VGND sg13g2_decap_4
X_10831_ _04843_ _04837_ _04839_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_450 VPWR VGND sg13g2_fill_2
X_13550_ VPWR _00101_ net88 VGND sg13g2_inv_1
XFILLER_41_921 VPWR VGND sg13g2_decap_8
XFILLER_16_63 VPWR VGND sg13g2_decap_8
XFILLER_16_74 VPWR VGND sg13g2_fill_1
X_10762_ _04774_ _04741_ VPWR VGND sg13g2_inv_2
XFILLER_25_483 VPWR VGND sg13g2_decap_8
X_12501_ VGND VPWR _03327_ net1951 _00957_ _06334_ sg13g2_a21oi_1
X_13481_ VPWR _00032_ net21 VGND sg13g2_inv_1
XFILLER_13_645 VPWR VGND sg13g2_decap_8
X_12432_ _06265_ _06277_ _06278_ VPWR VGND sg13g2_nor2b_1
XFILLER_40_475 VPWR VGND sg13g2_decap_4
XFILLER_8_126 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_decap_8
XFILLER_12_166 VPWR VGND sg13g2_decap_8
X_10693_ _04706_ _04704_ _04623_ VPWR VGND sg13g2_nand2_1
XFILLER_120_0 VPWR VGND sg13g2_decap_8
X_12363_ _06188_ _06208_ _06187_ _06209_ VPWR VGND sg13g2_nand3_1
XFILLER_5_822 VPWR VGND sg13g2_decap_8
X_12294_ _05974_ _05975_ _06137_ _06140_ VPWR VGND sg13g2_nand3_1
X_11314_ _01080_ _05269_ _05270_ VPWR VGND sg13g2_nand2_1
X_14102_ VPWR _00653_ net43 VGND sg13g2_inv_1
X_14033_ VPWR _00584_ net98 VGND sg13g2_inv_1
X_11245_ _02951_ _05194_ _05209_ VPWR VGND sg13g2_nor2_1
XFILLER_5_899 VPWR VGND sg13g2_decap_8
XFILLER_4_365 VPWR VGND sg13g2_decap_8
XFILLER_122_742 VPWR VGND sg13g2_decap_8
XFILLER_79_111 VPWR VGND sg13g2_decap_8
XFILLER_121_252 VPWR VGND sg13g2_decap_8
X_11176_ _05024_ _05144_ _05145_ VPWR VGND sg13g2_nor2_1
XFILLER_110_948 VPWR VGND sg13g2_decap_8
XFILLER_95_637 VPWR VGND sg13g2_decap_8
X_10127_ _04208_ VPWR _04209_ VGND _03611_ _04140_ sg13g2_o21ai_1
XFILLER_94_136 VPWR VGND sg13g2_decap_8
X_14935_ _00736_ VGND VPWR _01455_ acc_sub.exp_mant_logic0.a\[3\] clknet_leaf_56_clk
+ sg13g2_dfrbpq_2
X_10058_ _04017_ _04145_ _04146_ VPWR VGND sg13g2_nor2_1
XFILLER_36_715 VPWR VGND sg13g2_fill_2
XFILLER_36_704 VPWR VGND sg13g2_fill_1
XFILLER_91_865 VPWR VGND sg13g2_decap_4
XFILLER_91_832 VPWR VGND sg13g2_decap_4
XFILLER_35_225 VPWR VGND sg13g2_decap_4
XFILLER_17_940 VPWR VGND sg13g2_decap_8
X_14866_ _00667_ VGND VPWR _01390_ fp16_sum_pipe.seg_reg0.q\[28\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_1
X_13817_ VPWR _00368_ net77 VGND sg13g2_inv_1
X_14797_ _00598_ VGND VPWR _01321_ acc_sum.exp_mant_logic0.a\[10\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_13748_ VPWR _00299_ net123 VGND sg13g2_inv_1
XFILLER_31_420 VPWR VGND sg13g2_decap_8
XFILLER_32_943 VPWR VGND sg13g2_decap_8
XFILLER_31_453 VPWR VGND sg13g2_decap_4
X_13679_ VPWR _00230_ net120 VGND sg13g2_inv_1
XFILLER_31_497 VPWR VGND sg13g2_decap_8
XFILLER_117_569 VPWR VGND sg13g2_fill_1
XFILLER_117_558 VPWR VGND sg13g2_fill_2
X_09910_ _04004_ _04006_ _04007_ VPWR VGND sg13g2_nor2_1
XFILLER_99_965 VPWR VGND sg13g2_decap_8
XFILLER_113_753 VPWR VGND sg13g2_decap_8
X_09841_ net1803 _03949_ _03947_ _03952_ VPWR VGND _03951_ sg13g2_nand4_1
XFILLER_101_948 VPWR VGND sg13g2_decap_8
X_09772_ _03888_ _03827_ _03887_ VPWR VGND sg13g2_nand2_1
XFILLER_85_103 VPWR VGND sg13g2_decap_4
X_08723_ _02929_ net1819 acc_sum.seg_reg0.q\[24\] VPWR VGND sg13g2_nand2_1
XFILLER_39_542 VPWR VGND sg13g2_decap_8
XFILLER_85_169 VPWR VGND sg13g2_fill_2
XFILLER_82_821 VPWR VGND sg13g2_fill_1
X_08654_ _02874_ _02790_ _02873_ VPWR VGND sg13g2_xnor2_1
XFILLER_93_180 VPWR VGND sg13g2_fill_1
XFILLER_81_320 VPWR VGND sg13g2_decap_8
XFILLER_54_534 VPWR VGND sg13g2_decap_8
XFILLER_54_523 VPWR VGND sg13g2_fill_1
XFILLER_26_225 VPWR VGND sg13g2_decap_8
X_07605_ VPWR _01919_ _01918_ VGND sg13g2_inv_1
X_08585_ acc_sum.reg2en.q\[0\] VPWR _02808_ VGND _02807_ _02724_ sg13g2_o21ai_1
XFILLER_82_898 VPWR VGND sg13g2_decap_8
XFILLER_82_865 VPWR VGND sg13g2_decap_8
XFILLER_81_364 VPWR VGND sg13g2_decap_8
XFILLER_42_707 VPWR VGND sg13g2_decap_8
X_07536_ _01855_ _01844_ VPWR VGND sg13g2_inv_2
XFILLER_53_28 VPWR VGND sg13g2_decap_8
XFILLER_23_954 VPWR VGND sg13g2_decap_8
X_07467_ acc_sub.exp_mant_logic0.a\[14\] _01789_ _01790_ VPWR VGND sg13g2_nor2_1
X_09206_ fp16_res_pipe.reg2en.q\[0\] _03361_ VPWR VGND sg13g2_inv_4
X_07398_ _01740_ VPWR _01459_ VGND net1895 _01739_ sg13g2_o21ai_1
X_09137_ _03315_ VPWR _03316_ VGND _03165_ _03089_ sg13g2_o21ai_1
XFILLER_118_21 VPWR VGND sg13g2_decap_8
X_09068_ VGND VPWR _03252_ _03211_ _03253_ _03096_ sg13g2_a21oi_1
XFILLER_108_569 VPWR VGND sg13g2_decap_8
XFILLER_108_536 VPWR VGND sg13g2_fill_2
XFILLER_2_814 VPWR VGND sg13g2_decap_8
X_08019_ VPWR _02285_ _02284_ VGND sg13g2_inv_1
XFILLER_123_539 VPWR VGND sg13g2_decap_8
XFILLER_118_98 VPWR VGND sg13g2_decap_8
XFILLER_78_58 VPWR VGND sg13g2_decap_8
Xclkbuf_5_13__f_clk clknet_4_6_0_clk clknet_5_13__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_1_313 VPWR VGND sg13g2_fill_1
XFILLER_103_252 VPWR VGND sg13g2_fill_2
XFILLER_89_453 VPWR VGND sg13g2_decap_8
XFILLER_89_442 VPWR VGND sg13g2_fill_1
X_11030_ _05009_ _05008_ VPWR VGND sg13g2_inv_2
XFILLER_77_626 VPWR VGND sg13g2_decap_8
XFILLER_76_114 VPWR VGND sg13g2_decap_8
XFILLER_94_35 VPWR VGND sg13g2_fill_2
XFILLER_58_862 VPWR VGND sg13g2_decap_4
XFILLER_58_840 VPWR VGND sg13g2_decap_8
XFILLER_40_1013 VPWR VGND sg13g2_fill_1
XFILLER_73_821 VPWR VGND sg13g2_fill_1
XFILLER_64_309 VPWR VGND sg13g2_decap_8
X_12981_ VPWR _06749_ fpmul.seg_reg0.q\[20\] VGND sg13g2_inv_1
XFILLER_72_331 VPWR VGND sg13g2_decap_8
X_11932_ _05798_ VPWR _00990_ VGND net1879 _05797_ sg13g2_o21ai_1
X_14720_ _00521_ VGND VPWR _01248_ fp16_res_pipe.exp_mant_logic0.a\[7\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_2
XFILLER_73_876 VPWR VGND sg13g2_decap_8
X_14651_ _00452_ VGND VPWR _01179_ fp16_res_pipe.exp_mant_logic0.b\[4\] clknet_leaf_140_clk
+ sg13g2_dfrbpq_2
XFILLER_27_84 VPWR VGND sg13g2_decap_8
X_11863_ _05760_ _05759_ _05756_ VPWR VGND sg13g2_nand2b_1
X_13602_ VPWR _00153_ net121 VGND sg13g2_inv_1
XFILLER_72_397 VPWR VGND sg13g2_decap_8
XFILLER_60_537 VPWR VGND sg13g2_fill_1
X_10814_ VGND VPWR _04724_ _04808_ _04826_ _04825_ sg13g2_a21oi_1
XFILLER_32_206 VPWR VGND sg13g2_decap_8
XFILLER_32_217 VPWR VGND sg13g2_fill_2
XFILLER_41_751 VPWR VGND sg13g2_fill_2
XFILLER_41_740 VPWR VGND sg13g2_decap_8
X_14582_ _00383_ VGND VPWR _01114_ fp16_sum_pipe.exp_mant_logic0.b\[9\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_1
X_11794_ _05695_ _05608_ _05612_ _05696_ VPWR VGND sg13g2_a21o_1
XFILLER_14_965 VPWR VGND sg13g2_decap_8
X_13533_ VPWR _00084_ net85 VGND sg13g2_inv_1
XFILLER_41_795 VPWR VGND sg13g2_fill_1
X_10745_ _04758_ _04757_ net1771 VPWR VGND sg13g2_nand2_1
X_13464_ _07111_ VPWR _00772_ VGND _06937_ net1753 sg13g2_o21ai_1
XFILLER_40_294 VPWR VGND sg13g2_decap_8
X_10676_ VPWR _04689_ _04688_ VGND sg13g2_inv_1
XFILLER_127_834 VPWR VGND sg13g2_decap_8
X_13395_ _07074_ net1696 sipo.word\[1\] VPWR VGND sg13g2_nand2_1
X_12415_ _06051_ _06048_ _06261_ VPWR VGND sg13g2_and2_1
XFILLER_9_479 VPWR VGND sg13g2_decap_8
XFILLER_126_322 VPWR VGND sg13g2_decap_8
X_12346_ _06192_ net1858 net1868 VPWR VGND sg13g2_nand2_1
XFILLER_114_506 VPWR VGND sg13g2_decap_8
XFILLER_99_206 VPWR VGND sg13g2_decap_8
XFILLER_57_7 VPWR VGND sg13g2_decap_4
XFILLER_4_140 VPWR VGND sg13g2_decap_8
X_12277_ _05965_ _05971_ _06119_ _06123_ VPWR VGND sg13g2_nand3_1
X_14016_ VPWR _00567_ net75 VGND sg13g2_inv_1
XFILLER_4_77 VPWR VGND sg13g2_decap_8
X_11159_ _05128_ VPWR _01093_ VGND net1760 _05127_ sg13g2_o21ai_1
XFILLER_95_434 VPWR VGND sg13g2_fill_1
XFILLER_49_840 VPWR VGND sg13g2_decap_8
XFILLER_36_501 VPWR VGND sg13g2_fill_1
X_14918_ _00719_ VGND VPWR _01438_ acc_sub.seg_reg0.q\[28\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_82_139 VPWR VGND sg13g2_decap_4
XFILLER_64_887 VPWR VGND sg13g2_decap_4
XFILLER_63_342 VPWR VGND sg13g2_decap_8
XFILLER_51_504 VPWR VGND sg13g2_fill_1
X_14849_ _00650_ VGND VPWR _01373_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[0\] clknet_leaf_114_clk
+ sg13g2_dfrbpq_1
XFILLER_91_684 VPWR VGND sg13g2_decap_8
X_08370_ _02613_ _02611_ instr\[1\] _02612_ VPWR VGND sg13g2_and3_1
XFILLER_51_526 VPWR VGND sg13g2_decap_4
XFILLER_23_206 VPWR VGND sg13g2_decap_4
X_07321_ VPWR _01684_ _01563_ VGND sg13g2_inv_1
XFILLER_16_280 VPWR VGND sg13g2_fill_2
XFILLER_23_239 VPWR VGND sg13g2_decap_8
XFILLER_20_913 VPWR VGND sg13g2_decap_8
X_07252_ _01622_ net1783 acc_sub.add_renorm0.mantisa\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_83_0 VPWR VGND sg13g2_decap_8
XFILLER_31_272 VPWR VGND sg13g2_fill_2
X_07183_ acc_sub.op_sign_logic0.mantisa_a\[3\] _01554_ _01555_ VPWR VGND sg13g2_nor2_1
XFILLER_118_845 VPWR VGND sg13g2_decap_8
XFILLER_8_490 VPWR VGND sg13g2_decap_8
XFILLER_105_506 VPWR VGND sg13g2_decap_8
XFILLER_117_399 VPWR VGND sg13g2_fill_2
XFILLER_98_250 VPWR VGND sg13g2_decap_8
X_09824_ net1664 VPWR _03936_ VGND _03935_ _03925_ sg13g2_o21ai_1
XFILLER_59_626 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_87_979 VPWR VGND sg13g2_decap_8
XFILLER_86_434 VPWR VGND sg13g2_fill_2
X_09755_ _03857_ _03870_ _03871_ VPWR VGND sg13g2_nor2_2
XFILLER_104_45 VPWR VGND sg13g2_fill_1
XFILLER_55_810 VPWR VGND sg13g2_decap_4
X_09686_ _03802_ _03801_ acc_sum.add_renorm0.mantisa\[11\] VPWR VGND sg13g2_nand2_1
X_08706_ VPWR _02918_ acc_sum.add_renorm0.mantisa\[0\] VGND sg13g2_inv_1
XFILLER_27_534 VPWR VGND sg13g2_fill_1
X_08637_ _02837_ VPWR _02859_ VGND _02857_ _02858_ sg13g2_o21ai_1
XFILLER_70_802 VPWR VGND sg13g2_fill_1
XFILLER_55_887 VPWR VGND sg13g2_decap_8
XFILLER_81_172 VPWR VGND sg13g2_decap_8
XFILLER_70_846 VPWR VGND sg13g2_decap_8
X_08568_ _02788_ _02791_ _02792_ VPWR VGND sg13g2_nor2_1
Xfanout21 net23 net21 VPWR VGND sg13g2_buf_2
Xfanout10 net15 net10 VPWR VGND sg13g2_buf_2
XFILLER_120_77 VPWR VGND sg13g2_decap_8
X_07519_ _01840_ _01837_ _01821_ VPWR VGND sg13g2_nand2_1
X_08499_ acc_sum.op_sign_logic0.s_b acc_sum.op_sign_logic0.s_a _02724_ VPWR VGND sg13g2_xor2_1
Xfanout32 net34 net32 VPWR VGND sg13g2_buf_2
Xfanout54 net55 net54 VPWR VGND sg13g2_buf_2
Xfanout65 net66 net65 VPWR VGND sg13g2_buf_2
XFILLER_11_924 VPWR VGND sg13g2_decap_8
Xfanout43 net46 net43 VPWR VGND sg13g2_buf_2
XFILLER_23_762 VPWR VGND sg13g2_decap_8
Xfanout98 net100 net98 VPWR VGND sg13g2_buf_2
Xfanout87 net88 net87 VPWR VGND sg13g2_buf_2
Xfanout76 net93 net76 VPWR VGND sg13g2_buf_2
X_10530_ VGND VPWR net1670 _04506_ _04570_ net1737 sg13g2_a21oi_1
XFILLER_10_434 VPWR VGND sg13g2_decap_8
XFILLER_13_42 VPWR VGND sg13g2_decap_8
XFILLER_127_119 VPWR VGND sg13g2_decap_8
X_10461_ VGND VPWR _04508_ _04426_ _04509_ _04425_ sg13g2_a21oi_1
XFILLER_109_856 VPWR VGND sg13g2_decap_8
XFILLER_108_311 VPWR VGND sg13g2_fill_1
X_12200_ _06046_ _06043_ _06045_ VPWR VGND sg13g2_nand2_1
XFILLER_108_377 VPWR VGND sg13g2_decap_8
X_10392_ _04439_ _04441_ _04442_ VPWR VGND sg13g2_nor2_1
XFILLER_124_837 VPWR VGND sg13g2_decap_8
XFILLER_123_325 VPWR VGND sg13g2_decap_8
XFILLER_108_399 VPWR VGND sg13g2_fill_2
XFILLER_89_68 VPWR VGND sg13g2_decap_8
X_12131_ VGND VPWR _05974_ _05975_ _05977_ _05976_ sg13g2_a21oi_1
XFILLER_2_622 VPWR VGND sg13g2_decap_4
XFILLER_2_600 VPWR VGND sg13g2_decap_4
XFILLER_123_358 VPWR VGND sg13g2_decap_4
X_12062_ VPWR _05908_ _05907_ VGND sg13g2_inv_1
X_11013_ VPWR _04992_ acc_sum.seg_reg0.q\[29\] VGND sg13g2_inv_1
XFILLER_2_688 VPWR VGND sg13g2_fill_2
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_93_905 VPWR VGND sg13g2_decap_4
XFILLER_77_445 VPWR VGND sg13g2_decap_4
XFILLER_49_147 VPWR VGND sg13g2_decap_4
XFILLER_92_404 VPWR VGND sg13g2_decap_8
XFILLER_58_670 VPWR VGND sg13g2_fill_2
XFILLER_18_501 VPWR VGND sg13g2_fill_1
XFILLER_92_448 VPWR VGND sg13g2_decap_8
X_12964_ _06735_ _06734_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_46_843 VPWR VGND sg13g2_decap_8
XFILLER_18_523 VPWR VGND sg13g2_decap_8
X_14703_ _00504_ VGND VPWR _01231_ acc_sum.y\[6\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_46_854 VPWR VGND sg13g2_decap_4
X_11915_ VPWR _05787_ fpmul.seg_reg0.q\[41\] VGND sg13g2_inv_1
XFILLER_33_504 VPWR VGND sg13g2_decap_8
X_12895_ _00012_ net1731 net1702 _06671_ VPWR VGND sg13g2_nand3_1
XFILLER_73_695 VPWR VGND sg13g2_fill_1
XFILLER_73_673 VPWR VGND sg13g2_decap_8
XFILLER_45_397 VPWR VGND sg13g2_decap_4
XFILLER_45_386 VPWR VGND sg13g2_fill_2
XFILLER_33_515 VPWR VGND sg13g2_decap_8
XFILLER_33_526 VPWR VGND sg13g2_fill_2
XFILLER_61_868 VPWR VGND sg13g2_fill_1
XFILLER_61_857 VPWR VGND sg13g2_decap_4
X_14634_ _00435_ VGND VPWR _01166_ fp16_sum_pipe.add_renorm0.mantisa\[5\] clknet_leaf_108_clk
+ sg13g2_dfrbpq_2
X_11846_ _05635_ _05636_ _05742_ _05744_ VPWR VGND sg13g2_nand3_1
X_14565_ _00366_ VGND VPWR _01101_ acc_sum.seg_reg0.q\[28\] clknet_leaf_32_clk sg13g2_dfrbpq_1
X_11777_ fp16_sum_pipe.reg3en.q\[0\] _05679_ _05570_ _05680_ VPWR VGND sg13g2_nand3_1
X_13516_ VPWR _00067_ net89 VGND sg13g2_inv_1
XFILLER_14_795 VPWR VGND sg13g2_fill_1
X_10728_ _04741_ _04693_ _04740_ VPWR VGND sg13g2_nand2_2
XFILLER_118_119 VPWR VGND sg13g2_decap_8
X_14496_ _00297_ VGND VPWR _01032_ fpdiv.divider0.divisor\[7\] clknet_leaf_84_clk
+ sg13g2_dfrbpq_1
Xclkload13 clknet_5_27__leaf_clk clkload13/X VPWR VGND sg13g2_buf_8
Xclkload35 clknet_leaf_5_clk clkload35/X VPWR VGND sg13g2_buf_8
X_13447_ _07103_ net1754 sipo.shift_reg\[10\] VPWR VGND sg13g2_nand2_1
Xclkload24 VPWR clkload24/Y clknet_leaf_137_clk VGND sg13g2_inv_1
X_10659_ _04672_ fp16_res_pipe.add_renorm0.mantisa\[4\] _04641_ VPWR VGND sg13g2_xnor2_1
XFILLER_127_686 VPWR VGND sg13g2_decap_8
Xclkload68 clknet_leaf_27_clk clkload68/X VPWR VGND sg13g2_buf_8
Xclkload57 clkload57/Y clknet_leaf_94_clk VPWR VGND sg13g2_inv_8
X_13378_ _07065_ VPWR _00812_ VGND _06341_ net1694 sg13g2_o21ai_1
Xclkload46 clkload46/Y clknet_leaf_122_clk VPWR VGND sg13g2_inv_2
XFILLER_127_697 VPWR VGND sg13g2_fill_1
XFILLER_126_196 VPWR VGND sg13g2_decap_8
XFILLER_115_837 VPWR VGND sg13g2_decap_8
Xclkload79 clkload79/Y clknet_leaf_33_clk VPWR VGND sg13g2_inv_8
X_12329_ _06160_ _06167_ _06175_ VPWR VGND sg13g2_nor2_1
XFILLER_6_983 VPWR VGND sg13g2_decap_8
XFILLER_5_471 VPWR VGND sg13g2_decap_8
XFILLER_87_209 VPWR VGND sg13g2_decap_8
XFILLER_122_391 VPWR VGND sg13g2_fill_1
XFILLER_122_380 VPWR VGND sg13g2_decap_8
XFILLER_110_531 VPWR VGND sg13g2_decap_8
X_07870_ _02162_ net1888 acc_sub.x2\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_68_445 VPWR VGND sg13g2_fill_1
XFILLER_84_938 VPWR VGND sg13g2_decap_8
XFILLER_83_404 VPWR VGND sg13g2_decap_8
XFILLER_49_670 VPWR VGND sg13g2_decap_4
X_09540_ _03654_ _03655_ _03633_ _03657_ VPWR VGND sg13g2_nand3_1
XFILLER_110_1011 VPWR VGND sg13g2_fill_2
XFILLER_110_597 VPWR VGND sg13g2_fill_1
XFILLER_110_586 VPWR VGND sg13g2_fill_2
XFILLER_95_286 VPWR VGND sg13g2_decap_4
XFILLER_83_448 VPWR VGND sg13g2_decap_8
XFILLER_92_960 VPWR VGND sg13g2_decap_8
XFILLER_83_459 VPWR VGND sg13g2_fill_2
X_09471_ _03598_ VPWR _01251_ VGND net1914 _03597_ sg13g2_o21ai_1
XFILLER_36_353 VPWR VGND sg13g2_decap_8
X_08422_ VPWR _02656_ fpdiv.divider0.remainder_reg\[9\] VGND sg13g2_inv_1
XFILLER_64_673 VPWR VGND sg13g2_fill_1
XFILLER_24_515 VPWR VGND sg13g2_fill_1
XFILLER_91_492 VPWR VGND sg13g2_decap_8
XFILLER_52_857 VPWR VGND sg13g2_decap_8
X_08353_ instr\[11\] instr\[10\] instr\[9\] instr\[8\] _02596_ VPWR VGND sg13g2_nor4_1
XFILLER_51_367 VPWR VGND sg13g2_decap_8
X_07304_ net1744 _01608_ _01669_ _01670_ VPWR VGND sg13g2_nand3_1
X_08284_ _02531_ VPWR _02532_ VGND _02468_ _02345_ sg13g2_o21ai_1
XFILLER_32_570 VPWR VGND sg13g2_fill_1
X_07235_ _01606_ _01605_ _01536_ VPWR VGND sg13g2_nand2_1
Xclkload7 clknet_5_15__leaf_clk clkload7/X VPWR VGND sg13g2_buf_8
XFILLER_20_798 VPWR VGND sg13g2_decap_4
X_07166_ acc_sub.op_sign_logic0.mantisa_b\[4\] _01537_ _01538_ VPWR VGND sg13g2_nor2_1
XFILLER_106_804 VPWR VGND sg13g2_fill_2
XFILLER_4_909 VPWR VGND sg13g2_decap_8
XFILLER_118_697 VPWR VGND sg13g2_fill_1
XFILLER_59_16 VPWR VGND sg13g2_decap_8
XFILLER_117_196 VPWR VGND sg13g2_decap_8
XFILLER_59_49 VPWR VGND sg13g2_decap_8
XFILLER_114_881 VPWR VGND sg13g2_decap_8
XFILLER_101_531 VPWR VGND sg13g2_decap_4
XFILLER_87_765 VPWR VGND sg13g2_fill_1
XFILLER_59_456 VPWR VGND sg13g2_decap_8
XFILLER_115_77 VPWR VGND sg13g2_decap_8
X_09807_ _03920_ VPWR _01237_ VGND _03905_ _03919_ sg13g2_o21ai_1
XFILLER_75_927 VPWR VGND sg13g2_decap_8
XFILLER_74_415 VPWR VGND sg13g2_decap_8
XFILLER_19_309 VPWR VGND sg13g2_fill_1
X_07999_ _02186_ _02197_ _02238_ _02266_ VPWR VGND _02192_ sg13g2_nand4_1
X_09738_ _03854_ _03678_ _03849_ VPWR VGND sg13g2_nand2_1
XFILLER_74_426 VPWR VGND sg13g2_fill_2
XFILLER_90_919 VPWR VGND sg13g2_fill_2
XFILLER_83_960 VPWR VGND sg13g2_decap_8
XFILLER_55_662 VPWR VGND sg13g2_fill_1
XFILLER_43_802 VPWR VGND sg13g2_fill_1
XFILLER_39_191 VPWR VGND sg13g2_decap_4
XFILLER_28_854 VPWR VGND sg13g2_fill_1
XFILLER_55_695 VPWR VGND sg13g2_decap_4
XFILLER_54_172 VPWR VGND sg13g2_fill_1
XFILLER_70_632 VPWR VGND sg13g2_fill_2
X_12680_ _00937_ _06489_ _06492_ _06354_ _06488_ VPWR VGND sg13g2_a22oi_1
XFILLER_43_846 VPWR VGND sg13g2_decap_4
X_11700_ _05603_ VPWR _05604_ VGND _04587_ net1727 sg13g2_o21ai_1
X_11631_ _05535_ _05525_ _05531_ _05536_ VPWR VGND sg13g2_nor3_1
X_14350_ _00151_ VGND VPWR _00892_ fpmul.reg_p_out\[14\] clknet_leaf_92_clk sg13g2_dfrbpq_1
X_11562_ _05467_ _05428_ _05465_ _05459_ _05442_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_63 VPWR VGND sg13g2_decap_8
X_13301_ VGND VPWR net1678 _07012_ _00837_ _07013_ sg13g2_a21oi_1
X_10513_ net1848 fp16_sum_pipe.add_renorm0.mantisa\[5\] _04556_ VPWR VGND sg13g2_nor2_1
XFILLER_11_765 VPWR VGND sg13g2_decap_4
X_14281_ _00082_ VGND VPWR _00832_ fp16_res_pipe.x2\[14\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_11493_ VPWR _05398_ fp16_sum_pipe.add_renorm0.mantisa\[7\] VGND sg13g2_inv_1
X_13232_ _06953_ _06954_ _06955_ _06956_ _06957_ VPWR VGND sg13g2_nor4_1
X_10444_ _04493_ _04403_ _04492_ _04472_ net1736 VPWR VGND sg13g2_a22oi_1
XFILLER_40_84 VPWR VGND sg13g2_decap_8
X_10375_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[3\] _04424_ _04425_ VPWR VGND sg13g2_nor2_1
XFILLER_3_931 VPWR VGND sg13g2_decap_8
XFILLER_123_133 VPWR VGND sg13g2_decap_8
X_12114_ _05960_ _05900_ _05959_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_430 VPWR VGND sg13g2_decap_8
X_13094_ _06855_ _06854_ _06805_ VPWR VGND sg13g2_nand2_1
X_12045_ _05891_ net1860 VPWR VGND sg13g2_inv_2
XFILLER_120_862 VPWR VGND sg13g2_decap_8
XFILLER_78_798 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_19_832 VPWR VGND sg13g2_decap_8
XFILLER_92_245 VPWR VGND sg13g2_fill_1
XFILLER_81_919 VPWR VGND sg13g2_fill_1
XFILLER_74_960 VPWR VGND sg13g2_decap_8
XFILLER_46_640 VPWR VGND sg13g2_fill_1
X_13996_ VPWR _00547_ net10 VGND sg13g2_inv_1
XFILLER_80_429 VPWR VGND sg13g2_decap_8
X_12947_ _06718_ _06717_ fp16_sum_pipe.reg1en.d\[0\] _06719_ VPWR VGND sg13g2_a21o_2
XFILLER_45_161 VPWR VGND sg13g2_decap_8
XFILLER_34_813 VPWR VGND sg13g2_decap_8
XFILLER_18_364 VPWR VGND sg13g2_decap_8
XFILLER_18_375 VPWR VGND sg13g2_fill_2
XFILLER_19_887 VPWR VGND sg13g2_decap_8
X_12878_ _06656_ _06655_ fpmul.reg1en.d\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_60_120 VPWR VGND sg13g2_decap_8
X_14617_ _00418_ VGND VPWR _01149_ fp16_sum_pipe.exp_mant_logic0.a\[12\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_2
X_11829_ _05729_ _05719_ _05728_ VPWR VGND sg13g2_nand2_1
XFILLER_21_507 VPWR VGND sg13g2_decap_8
XFILLER_61_698 VPWR VGND sg13g2_fill_2
X_14548_ _00349_ VGND VPWR _01084_ acc_sum.op_sign_logic0.mantisa_a\[0\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
XFILLER_14_1007 VPWR VGND sg13g2_decap_8
Xclkload113 clkload113/Y clknet_leaf_71_clk VPWR VGND sg13g2_inv_8
Xclkload102 clknet_leaf_76_clk clkload102/Y VPWR VGND sg13g2_inv_4
X_14479_ _00280_ VGND VPWR _01017_ add_result\[4\] clknet_leaf_107_clk sg13g2_dfrbpq_2
XFILLER_60_2 VPWR VGND sg13g2_fill_1
Xplace1903 net1902 net1903 VPWR VGND sg13g2_buf_2
Xplace1936 net1935 net1936 VPWR VGND sg13g2_buf_2
Xplace1914 net1913 net1914 VPWR VGND sg13g2_buf_2
Xplace1925 net1924 net1925 VPWR VGND sg13g2_buf_2
XFILLER_114_133 VPWR VGND sg13g2_decap_8
Xplace1947 net1946 net1947 VPWR VGND sg13g2_buf_2
Xplace1958 fpmul.reg1en.d\[0\] net1958 VPWR VGND sg13g2_buf_2
XFILLER_46_0 VPWR VGND sg13g2_decap_8
XFILLER_5_290 VPWR VGND sg13g2_decap_8
X_08971_ VGND VPWR _03156_ _03157_ _03155_ net1699 sg13g2_a21oi_2
XFILLER_88_529 VPWR VGND sg13g2_fill_1
XFILLER_68_231 VPWR VGND sg13g2_decap_4
X_07922_ _02197_ fp16_sum_pipe.exp_mant_logic0.a\[12\] VPWR VGND sg13g2_inv_2
XFILLER_111_873 VPWR VGND sg13g2_decap_8
X_07853_ _02148_ _02147_ net1640 VPWR VGND sg13g2_nand2_1
XFILLER_68_264 VPWR VGND sg13g2_decap_8
XFILLER_83_201 VPWR VGND sg13g2_decap_8
XFILLER_56_448 VPWR VGND sg13g2_decap_8
XFILLER_56_437 VPWR VGND sg13g2_fill_1
X_07784_ _02082_ _02083_ _02081_ _02084_ VPWR VGND sg13g2_nand3_1
XFILLER_84_779 VPWR VGND sg13g2_decap_8
XFILLER_25_802 VPWR VGND sg13g2_fill_1
X_09523_ _03640_ _03639_ _03625_ VPWR VGND sg13g2_nand2_2
XFILLER_25_835 VPWR VGND sg13g2_fill_1
XFILLER_101_13 VPWR VGND sg13g2_decap_8
XFILLER_24_345 VPWR VGND sg13g2_decap_8
X_09454_ fp16_res_pipe.add_renorm0.exp\[0\] fp16_res_pipe.seg_reg0.q\[22\] net1833
+ _01257_ VPWR VGND sg13g2_mux2_1
X_08405_ _02640_ _02633_ _02641_ VPWR VGND sg13g2_and2_1
XFILLER_40_805 VPWR VGND sg13g2_decap_8
X_09385_ _03533_ _03388_ _03470_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_378 VPWR VGND sg13g2_fill_2
X_08336_ _02563_ _02566_ _02569_ _02580_ _02581_ VPWR VGND sg13g2_nor4_1
XFILLER_61_28 VPWR VGND sg13g2_decap_4
XFILLER_33_890 VPWR VGND sg13g2_decap_8
XFILLER_124_7 VPWR VGND sg13g2_decap_8
XFILLER_119_940 VPWR VGND sg13g2_decap_8
X_08267_ _01366_ _02515_ _02516_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_140_clk clknet_5_0__leaf_clk clknet_leaf_140_clk VPWR VGND sg13g2_buf_8
X_07218_ _01580_ _01589_ _01590_ VPWR VGND _01502_ sg13g2_nand3b_1
X_08198_ _02455_ net1639 _02454_ VPWR VGND sg13g2_nand2_1
X_07149_ _01518_ _01520_ _01521_ VPWR VGND sg13g2_nor2_2
XFILLER_10_21 VPWR VGND sg13g2_decap_8
XFILLER_126_21 VPWR VGND sg13g2_decap_8
XFILLER_106_667 VPWR VGND sg13g2_decap_4
XFILLER_3_238 VPWR VGND sg13g2_decap_4
XFILLER_0_912 VPWR VGND sg13g2_decap_8
X_10160_ _04241_ _04240_ net1637 VPWR VGND sg13g2_nand2_1
XFILLER_126_98 VPWR VGND sg13g2_decap_8
XFILLER_121_659 VPWR VGND sg13g2_fill_1
XFILLER_105_199 VPWR VGND sg13g2_decap_8
XFILLER_86_47 VPWR VGND sg13g2_fill_2
XFILLER_10_98 VPWR VGND sg13g2_decap_8
XFILLER_120_147 VPWR VGND sg13g2_decap_8
XFILLER_87_562 VPWR VGND sg13g2_decap_8
XFILLER_0_989 VPWR VGND sg13g2_decap_8
XFILLER_74_223 VPWR VGND sg13g2_decap_8
XFILLER_19_63 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_fill_1
XFILLER_19_106 VPWR VGND sg13g2_decap_8
X_13850_ VPWR _00401_ net29 VGND sg13g2_inv_1
X_13781_ VPWR _00332_ net126 VGND sg13g2_inv_1
XFILLER_90_749 VPWR VGND sg13g2_fill_2
XFILLER_76_1012 VPWR VGND sg13g2_fill_2
XFILLER_74_278 VPWR VGND sg13g2_decap_8
X_12801_ _06585_ _06581_ _06584_ _06371_ net1941 VPWR VGND sg13g2_a22oi_1
XFILLER_27_161 VPWR VGND sg13g2_fill_2
X_10993_ _04982_ VPWR _01113_ VGND net1932 _02227_ sg13g2_o21ai_1
X_12732_ _06535_ VPWR _00928_ VGND _06533_ _02648_ sg13g2_o21ai_1
XFILLER_71_963 VPWR VGND sg13g2_fill_2
XFILLER_71_952 VPWR VGND sg13g2_decap_8
XFILLER_71_930 VPWR VGND sg13g2_decap_4
XFILLER_16_868 VPWR VGND sg13g2_decap_8
XFILLER_35_84 VPWR VGND sg13g2_decap_8
XFILLER_31_805 VPWR VGND sg13g2_fill_2
XFILLER_31_827 VPWR VGND sg13g2_decap_8
X_12663_ VGND VPWR _06354_ _06479_ _06360_ _06478_ sg13g2_a21oi_2
X_14402_ _00203_ VGND VPWR _00941_ div_result\[15\] clknet_leaf_90_clk sg13g2_dfrbpq_1
XFILLER_24_890 VPWR VGND sg13g2_decap_8
X_12594_ _06410_ fpdiv.reg_a_out\[13\] fpdiv.reg_b_out\[13\] VPWR VGND sg13g2_xnor2_1
X_11614_ VGND VPWR net1840 _05409_ _05519_ _05518_ sg13g2_a21oi_1
X_14333_ _00134_ VGND VPWR _00875_ piso.tx_bit_counter\[2\] clknet_leaf_57_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_131_clk clknet_5_3__leaf_clk clknet_leaf_131_clk VPWR VGND sg13g2_buf_8
XFILLER_11_573 VPWR VGND sg13g2_fill_2
X_11545_ _05450_ _05444_ _05449_ VPWR VGND sg13g2_nand2_1
X_11476_ _05390_ fp16_res_pipe.x2\[8\] net1942 VPWR VGND sg13g2_nand2_1
X_14264_ _00065_ VGND VPWR _00815_ acc_sub.x2\[13\] clknet_leaf_127_clk sg13g2_dfrbpq_2
XFILLER_125_921 VPWR VGND sg13g2_decap_8
X_13215_ VGND VPWR _06899_ _06880_ _06944_ sipo.bit_counter\[3\] sg13g2_a21oi_1
X_10427_ _04476_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[1\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[1\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_98_816 VPWR VGND sg13g2_fill_1
X_14195_ VPWR _00746_ net114 VGND sg13g2_inv_1
XFILLER_125_998 VPWR VGND sg13g2_decap_8
X_13146_ VGND VPWR piso.tx_bit_counter\[0\] _06882_ _00873_ _06894_ sg13g2_a21oi_1
X_10358_ _04405_ _04407_ _04408_ VPWR VGND sg13g2_nor2_2
X_13077_ VGND VPWR _06813_ _06757_ _06843_ _06835_ sg13g2_a21oi_1
X_10289_ _04358_ _04357_ net1636 VPWR VGND sg13g2_nand2_1
X_12028_ _05875_ VPWR _00971_ VGND net1873 _05873_ sg13g2_o21ai_1
XFILLER_2_293 VPWR VGND sg13g2_decap_4
XFILLER_66_757 VPWR VGND sg13g2_fill_1
XFILLER_54_908 VPWR VGND sg13g2_decap_8
XFILLER_38_448 VPWR VGND sg13g2_fill_2
XFILLER_20_1011 VPWR VGND sg13g2_fill_2
XFILLER_81_716 VPWR VGND sg13g2_decap_8
X_13979_ VPWR _00530_ net12 VGND sg13g2_inv_1
XFILLER_80_226 VPWR VGND sg13g2_fill_1
XFILLER_33_120 VPWR VGND sg13g2_decap_4
XFILLER_90_1009 VPWR VGND sg13g2_decap_4
XFILLER_34_687 VPWR VGND sg13g2_decap_8
XFILLER_61_495 VPWR VGND sg13g2_decap_8
XFILLER_119_203 VPWR VGND sg13g2_decap_8
X_09170_ _03336_ VPWR _01290_ VGND net1904 _03335_ sg13g2_o21ai_1
Xclkbuf_leaf_122_clk clknet_5_9__leaf_clk clknet_leaf_122_clk VPWR VGND sg13g2_buf_8
X_08121_ _02260_ net1648 _02383_ VPWR VGND sg13g2_nor2_1
XFILLER_30_871 VPWR VGND sg13g2_fill_1
X_08052_ _02318_ _02214_ _02317_ VPWR VGND sg13g2_xnor2_1
Xplace1711 _02578_ net1711 VPWR VGND sg13g2_buf_1
Xplace1700 _06837_ net1700 VPWR VGND sg13g2_buf_2
XFILLER_127_280 VPWR VGND sg13g2_decap_8
Xplace1744 _01496_ net1744 VPWR VGND sg13g2_buf_2
XFILLER_116_954 VPWR VGND sg13g2_decap_8
Xplace1733 net1732 net1733 VPWR VGND sg13g2_buf_2
Xplace1722 _07076_ net1722 VPWR VGND sg13g2_buf_2
XFILLER_103_626 VPWR VGND sg13g2_fill_2
Xplace1755 _06750_ net1755 VPWR VGND sg13g2_buf_2
Xplace1766 _03988_ net1766 VPWR VGND sg13g2_buf_1
Xplace1777 net1774 net1777 VPWR VGND sg13g2_buf_1
XFILLER_0_219 VPWR VGND sg13g2_fill_1
Xplace1788 acc_sub.add_renorm0.mantisa\[11\] net1788 VPWR VGND sg13g2_buf_2
X_08954_ _01717_ _03139_ _03140_ VPWR VGND sg13g2_nor2_1
Xplace1799 net1797 net1799 VPWR VGND sg13g2_buf_1
XFILLER_103_659 VPWR VGND sg13g2_decap_4
XFILLER_102_158 VPWR VGND sg13g2_decap_8
X_08885_ _03060_ VPWR _03072_ VGND _03062_ _03068_ sg13g2_o21ai_1
XFILLER_111_670 VPWR VGND sg13g2_decap_8
XFILLER_84_510 VPWR VGND sg13g2_decap_4
XFILLER_69_595 VPWR VGND sg13g2_decap_8
XFILLER_57_724 VPWR VGND sg13g2_decap_8
XFILLER_56_28 VPWR VGND sg13g2_fill_2
X_07836_ _02131_ VPWR _02132_ VGND _02130_ _01979_ sg13g2_o21ai_1
XFILLER_56_245 VPWR VGND sg13g2_decap_8
XFILLER_56_234 VPWR VGND sg13g2_decap_8
XFILLER_45_908 VPWR VGND sg13g2_fill_1
X_07767_ _02069_ net1685 net1795 VPWR VGND sg13g2_nand2_1
XFILLER_84_576 VPWR VGND sg13g2_decap_8
XFILLER_56_267 VPWR VGND sg13g2_decap_8
XFILLER_112_56 VPWR VGND sg13g2_decap_8
X_09506_ acc_sum.add_renorm0.mantisa\[5\] acc_sum.add_renorm0.mantisa\[4\] _03622_
+ _03623_ VPWR VGND sg13g2_nand3_1
XFILLER_25_643 VPWR VGND sg13g2_fill_1
X_07698_ _02005_ net1660 _02006_ VPWR VGND sg13g2_nor2_2
XFILLER_53_974 VPWR VGND sg13g2_decap_8
X_09437_ _03577_ net1834 fp16_res_pipe.seg_reg0.q\[28\] VPWR VGND sg13g2_nand2_1
XFILLER_12_304 VPWR VGND sg13g2_fill_1
XFILLER_13_849 VPWR VGND sg13g2_decap_8
XFILLER_25_698 VPWR VGND sg13g2_decap_8
XFILLER_40_679 VPWR VGND sg13g2_decap_8
X_09368_ _03501_ _03518_ VPWR VGND sg13g2_inv_4
X_08319_ state\[1\] state\[0\] _02564_ VPWR VGND sg13g2_nor2_1
X_09299_ VGND VPWR _03445_ _03453_ _03452_ _03440_ sg13g2_a21oi_2
XFILLER_21_882 VPWR VGND sg13g2_decap_8
X_11330_ _05285_ _05280_ _05284_ VPWR VGND sg13g2_nand2_1
XFILLER_20_392 VPWR VGND sg13g2_decap_8
XFILLER_126_729 VPWR VGND sg13g2_decap_8
XFILLER_125_217 VPWR VGND sg13g2_decap_8
XFILLER_4_525 VPWR VGND sg13g2_decap_8
XFILLER_21_42 VPWR VGND sg13g2_decap_8
XFILLER_107_943 VPWR VGND sg13g2_decap_8
X_11261_ _05223_ VPWR _05224_ VGND _02963_ _05222_ sg13g2_o21ai_1
XFILLER_122_924 VPWR VGND sg13g2_decap_8
X_13000_ _06767_ VPWR _06768_ VGND net1755 fpmul.seg_reg0.q\[14\] sg13g2_o21ai_1
X_10212_ _04287_ fp16_res_pipe.exp_mant_logic0.b\[4\] net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[7\]
+ net1763 VPWR VGND sg13g2_a22oi_1
XFILLER_97_68 VPWR VGND sg13g2_decap_4
X_10143_ _04224_ _04135_ VPWR VGND sg13g2_inv_2
XFILLER_0_764 VPWR VGND sg13g2_decap_8
X_14951_ _00752_ VGND VPWR _01471_ acc_sub.add_renorm0.exp\[3\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_94_329 VPWR VGND sg13g2_fill_1
XFILLER_48_724 VPWR VGND sg13g2_decap_8
XFILLER_0_786 VPWR VGND sg13g2_decap_8
X_10074_ _04159_ _04160_ _04155_ _04161_ VPWR VGND sg13g2_nand3_1
X_14882_ _00683_ VGND VPWR _01402_ acc_sub.exp_mant_logic0.b\[8\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_2
X_13902_ VPWR _00453_ net11 VGND sg13g2_inv_1
XFILLER_90_513 VPWR VGND sg13g2_fill_2
X_13833_ VPWR _00384_ net56 VGND sg13g2_inv_1
XFILLER_35_407 VPWR VGND sg13g2_decap_8
X_13764_ VPWR _00315_ net117 VGND sg13g2_inv_1
XFILLER_71_771 VPWR VGND sg13g2_fill_2
X_10976_ fp16_res_pipe.y\[1\] _04708_ net1835 _01122_ VPWR VGND sg13g2_mux2_1
XFILLER_43_462 VPWR VGND sg13g2_decap_8
XFILLER_15_131 VPWR VGND sg13g2_fill_1
XFILLER_16_665 VPWR VGND sg13g2_fill_2
X_12715_ _06521_ _06504_ _06423_ VPWR VGND sg13g2_nand2_1
X_13695_ VPWR _00246_ net70 VGND sg13g2_inv_1
XFILLER_15_175 VPWR VGND sg13g2_decap_8
XFILLER_31_624 VPWR VGND sg13g2_decap_8
XFILLER_87_7 VPWR VGND sg13g2_fill_1
X_12646_ _06462_ _06461_ _06419_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_145 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_104_clk clknet_5_14__leaf_clk clknet_leaf_104_clk VPWR VGND sg13g2_buf_8
XFILLER_117_718 VPWR VGND sg13g2_decap_8
X_12577_ _06391_ _06390_ _06393_ VPWR VGND sg13g2_and2_1
X_14316_ _00117_ VGND VPWR _00859_ sipo.word\[4\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_8_853 VPWR VGND sg13g2_decap_8
XFILLER_7_330 VPWR VGND sg13g2_fill_1
XFILLER_7_77 VPWR VGND sg13g2_decap_8
X_11528_ VPWR _05433_ _05426_ VGND sg13g2_inv_1
XFILLER_109_291 VPWR VGND sg13g2_decap_4
X_11459_ _05382_ acc_sub.x2\[1\] VPWR VGND sg13g2_inv_2
X_14247_ _00048_ VGND VPWR _00798_ instr\[12\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_98_613 VPWR VGND sg13g2_decap_8
X_14178_ VPWR _00729_ net127 VGND sg13g2_inv_1
XFILLER_125_795 VPWR VGND sg13g2_decap_8
XFILLER_124_294 VPWR VGND sg13g2_decap_8
XFILLER_113_935 VPWR VGND sg13g2_decap_8
XFILLER_112_423 VPWR VGND sg13g2_decap_8
X_13129_ VGND VPWR _06882_ _06881_ _06556_ sg13g2_or2_1
XFILLER_3_580 VPWR VGND sg13g2_decap_8
XFILLER_100_618 VPWR VGND sg13g2_fill_1
XFILLER_97_167 VPWR VGND sg13g2_fill_1
XFILLER_66_521 VPWR VGND sg13g2_decap_8
X_08670_ net1818 acc_sum.add_renorm0.mantisa\[6\] _02888_ VPWR VGND sg13g2_nor2_1
XFILLER_66_532 VPWR VGND sg13g2_fill_1
XFILLER_39_768 VPWR VGND sg13g2_decap_8
X_07621_ _01905_ _01934_ _01935_ VPWR VGND sg13g2_nor2b_2
XFILLER_66_576 VPWR VGND sg13g2_fill_2
XFILLER_53_204 VPWR VGND sg13g2_decap_8
X_07552_ _01747_ _01749_ _01741_ _01867_ VPWR VGND _01753_ sg13g2_nand4_1
XFILLER_19_481 VPWR VGND sg13g2_decap_8
XFILLER_35_974 VPWR VGND sg13g2_decap_8
X_07483_ _01803_ _01805_ _01806_ VPWR VGND sg13g2_nor2_1
XFILLER_50_922 VPWR VGND sg13g2_decap_8
XFILLER_22_613 VPWR VGND sg13g2_decap_4
XFILLER_22_624 VPWR VGND sg13g2_decap_4
X_09222_ _03376_ _03374_ _03375_ VPWR VGND sg13g2_nand2_2
X_09153_ _03325_ VPWR _01296_ VGND net1773 _03125_ sg13g2_o21ai_1
X_09084_ VGND VPWR _03251_ _03267_ _03268_ _03096_ sg13g2_a21oi_1
X_08035_ _02286_ _02245_ _02301_ VPWR VGND sg13g2_nor2_1
XFILLER_116_751 VPWR VGND sg13g2_decap_8
XFILLER_101_9 VPWR VGND sg13g2_fill_1
XFILLER_89_613 VPWR VGND sg13g2_decap_4
XFILLER_1_506 VPWR VGND sg13g2_decap_8
XFILLER_104_957 VPWR VGND sg13g2_decap_8
XFILLER_88_112 VPWR VGND sg13g2_decap_4
X_09986_ fp16_res_pipe.reg1en.q\[0\] _04073_ _04047_ _04075_ VPWR VGND sg13g2_nand3_1
X_08937_ acc_sub.seg_reg1.q\[21\] _03032_ _03123_ _03124_ VPWR VGND sg13g2_nor3_1
XFILLER_67_49 VPWR VGND sg13g2_decap_4
X_08868_ _01490_ _02979_ _03055_ VPWR VGND sg13g2_nor2_1
XFILLER_123_77 VPWR VGND sg13g2_decap_8
X_07819_ _02116_ net1646 acc_sub.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_84_373 VPWR VGND sg13g2_decap_4
XFILLER_57_587 VPWR VGND sg13g2_fill_2
XFILLER_17_418 VPWR VGND sg13g2_decap_8
X_08799_ VGND VPWR _01700_ _01707_ _02986_ _02985_ sg13g2_a21oi_1
XFILLER_84_384 VPWR VGND sg13g2_decap_8
XFILLER_83_59 VPWR VGND sg13g2_fill_2
XFILLER_72_535 VPWR VGND sg13g2_decap_4
XFILLER_44_215 VPWR VGND sg13g2_fill_2
XFILLER_60_708 VPWR VGND sg13g2_decap_8
XFILLER_16_42 VPWR VGND sg13g2_decap_8
X_10830_ VPWR _04842_ _04841_ VGND sg13g2_inv_1
X_10761_ _04773_ VPWR _01136_ VGND _03367_ _04771_ sg13g2_o21ai_1
XFILLER_26_996 VPWR VGND sg13g2_decap_8
X_12500_ fpmul.reg_a_out\[15\] net1951 _06334_ VPWR VGND sg13g2_nor2_1
XFILLER_52_292 VPWR VGND sg13g2_decap_4
X_13480_ VPWR _00031_ net21 VGND sg13g2_inv_1
XFILLER_9_606 VPWR VGND sg13g2_decap_8
XFILLER_12_112 VPWR VGND sg13g2_fill_2
X_10692_ _04623_ _04704_ _04705_ VPWR VGND sg13g2_nor2_1
X_12431_ _06277_ _06275_ _06276_ VPWR VGND sg13g2_xnor2_1
XFILLER_8_105 VPWR VGND sg13g2_decap_8
XFILLER_9_639 VPWR VGND sg13g2_decap_4
XFILLER_32_63 VPWR VGND sg13g2_decap_8
X_12362_ VPWR _06208_ _06207_ VGND sg13g2_inv_1
XFILLER_113_0 VPWR VGND sg13g2_decap_8
X_12293_ _06139_ _06138_ _05975_ VPWR VGND sg13g2_nand2b_1
X_11313_ _05270_ acc_sum.exp_mant_logic0.b\[4\] net1681 acc_sum.op_sign_logic0.mantisa_b\[7\]
+ net1762 VPWR VGND sg13g2_a22oi_1
X_14101_ VPWR _00652_ net42 VGND sg13g2_inv_1
XFILLER_10_1010 VPWR VGND sg13g2_decap_4
XFILLER_113_209 VPWR VGND sg13g2_decap_8
X_14032_ VPWR _00583_ net98 VGND sg13g2_inv_1
X_11244_ _05208_ _05161_ acc_sum.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_5_878 VPWR VGND sg13g2_decap_8
XFILLER_4_344 VPWR VGND sg13g2_decap_8
XFILLER_122_721 VPWR VGND sg13g2_decap_8
XFILLER_106_272 VPWR VGND sg13g2_fill_1
XFILLER_106_261 VPWR VGND sg13g2_decap_8
XFILLER_121_231 VPWR VGND sg13g2_decap_8
XFILLER_79_156 VPWR VGND sg13g2_decap_8
X_11175_ _05144_ _05131_ VPWR VGND sg13g2_inv_2
XFILLER_67_307 VPWR VGND sg13g2_fill_1
XFILLER_122_798 VPWR VGND sg13g2_decap_8
XFILLER_110_927 VPWR VGND sg13g2_decap_8
XFILLER_94_115 VPWR VGND sg13g2_decap_8
XFILLER_79_167 VPWR VGND sg13g2_fill_1
X_10126_ _04208_ net1642 net1828 VPWR VGND sg13g2_nand2_1
X_14934_ _00735_ VGND VPWR _01454_ acc_sub.exp_mant_logic0.a\[2\] clknet_leaf_56_clk
+ sg13g2_dfrbpq_2
X_10057_ VPWR _04145_ _04128_ VGND sg13g2_inv_1
XFILLER_75_340 VPWR VGND sg13g2_fill_2
XFILLER_63_502 VPWR VGND sg13g2_fill_2
X_14865_ _00666_ VGND VPWR _01389_ fp16_sum_pipe.seg_reg0.q\[27\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_1
X_13816_ VPWR _00367_ net77 VGND sg13g2_inv_1
X_14796_ _00597_ VGND VPWR _01320_ acc_sum.exp_mant_logic0.a\[9\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_63_579 VPWR VGND sg13g2_decap_4
XFILLER_90_376 VPWR VGND sg13g2_fill_1
X_13747_ VPWR _00298_ net117 VGND sg13g2_inv_1
XFILLER_44_782 VPWR VGND sg13g2_decap_4
XFILLER_17_996 VPWR VGND sg13g2_decap_8
X_10959_ _04964_ _04739_ _04842_ VPWR VGND sg13g2_nand2_1
XFILLER_32_922 VPWR VGND sg13g2_decap_8
X_13678_ VPWR _00229_ net120 VGND sg13g2_inv_1
XFILLER_31_476 VPWR VGND sg13g2_decap_8
XFILLER_32_999 VPWR VGND sg13g2_decap_8
X_12629_ VPWR _06445_ _06444_ VGND sg13g2_inv_1
XFILLER_89_1000 VPWR VGND sg13g2_decap_8
XFILLER_117_504 VPWR VGND sg13g2_decap_8
XFILLER_99_944 VPWR VGND sg13g2_decap_8
X_09840_ _03663_ _03950_ _03951_ VPWR VGND _03879_ sg13g2_nand3b_1
X_09771_ _03887_ _03869_ _03886_ VPWR VGND sg13g2_nand2_1
XFILLER_101_927 VPWR VGND sg13g2_decap_8
XFILLER_39_510 VPWR VGND sg13g2_decap_8
X_08722_ VPWR _02928_ acc_sum.add_renorm0.exp\[2\] VGND sg13g2_inv_1
XFILLER_79_690 VPWR VGND sg13g2_fill_2
XFILLER_96_1004 VPWR VGND sg13g2_decap_8
XFILLER_67_896 VPWR VGND sg13g2_fill_1
XFILLER_67_863 VPWR VGND sg13g2_decap_8
XFILLER_26_204 VPWR VGND sg13g2_decap_8
X_08653_ VGND VPWR _02871_ _02872_ _02873_ _02834_ sg13g2_a21oi_1
XFILLER_66_395 VPWR VGND sg13g2_decap_8
XFILLER_66_373 VPWR VGND sg13g2_fill_2
X_07604_ _01918_ _01806_ _01917_ VPWR VGND sg13g2_xnor2_1
X_08584_ _02807_ acc_sum.op_sign_logic0.mantisa_a\[10\] acc_sum.op_sign_logic0.mantisa_b\[10\]
+ VPWR VGND sg13g2_nand2_1
X_07535_ _01853_ _01854_ _01852_ _01436_ VPWR VGND sg13g2_nand3_1
XFILLER_41_207 VPWR VGND sg13g2_fill_1
XFILLER_35_793 VPWR VGND sg13g2_fill_2
XFILLER_35_782 VPWR VGND sg13g2_decap_8
XFILLER_23_933 VPWR VGND sg13g2_decap_8
X_07466_ VPWR _01789_ acc_sub.exp_mant_logic0.b\[14\] VGND sg13g2_inv_1
XFILLER_50_785 VPWR VGND sg13g2_decap_8
XFILLER_10_616 VPWR VGND sg13g2_fill_2
XFILLER_22_476 VPWR VGND sg13g2_decap_8
XFILLER_120_1002 VPWR VGND sg13g2_decap_8
X_07397_ _01740_ net1893 acc\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_120_1013 VPWR VGND sg13g2_fill_1
X_09136_ VGND VPWR _03101_ _03165_ _03315_ net1785 sg13g2_a21oi_1
XFILLER_5_119 VPWR VGND sg13g2_decap_8
X_09067_ _03252_ _03251_ _03153_ VPWR VGND sg13g2_nand2_1
X_08018_ VGND VPWR _02283_ _02235_ _02284_ _02195_ sg13g2_a21oi_1
XFILLER_118_77 VPWR VGND sg13g2_decap_8
XFILLER_116_570 VPWR VGND sg13g2_decap_8
XFILLER_89_432 VPWR VGND sg13g2_fill_1
XFILLER_1_303 VPWR VGND sg13g2_fill_2
XFILLER_104_743 VPWR VGND sg13g2_decap_8
XFILLER_103_275 VPWR VGND sg13g2_fill_2
XFILLER_77_638 VPWR VGND sg13g2_fill_1
X_09969_ _04061_ VPWR _01216_ VGND _04018_ _04054_ sg13g2_o21ai_1
XFILLER_94_14 VPWR VGND sg13g2_decap_8
XFILLER_76_126 VPWR VGND sg13g2_decap_8
X_12980_ VPWR _06748_ fpmul.seg_reg0.q\[22\] VGND sg13g2_inv_1
XFILLER_100_993 VPWR VGND sg13g2_decap_8
XFILLER_91_129 VPWR VGND sg13g2_decap_8
XFILLER_72_310 VPWR VGND sg13g2_decap_8
X_11931_ _05798_ net1879 fpmul.reg_b_out\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_45_513 VPWR VGND sg13g2_decap_8
XFILLER_27_63 VPWR VGND sg13g2_decap_8
X_14650_ _00451_ VGND VPWR _01178_ fp16_res_pipe.exp_mant_logic0.b\[3\] clknet_leaf_140_clk
+ sg13g2_dfrbpq_2
X_11862_ _05758_ VPWR _05759_ VGND _05636_ _05489_ sg13g2_o21ai_1
XFILLER_72_387 VPWR VGND sg13g2_fill_1
X_13601_ VPWR _00152_ net108 VGND sg13g2_inv_1
X_14581_ _00382_ VGND VPWR _01113_ fp16_sum_pipe.exp_mant_logic0.b\[8\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_2
X_10813_ _04822_ _04824_ _04825_ VPWR VGND sg13g2_and2_1
X_13532_ VPWR _00083_ net37 VGND sg13g2_inv_1
X_11793_ _05695_ _05601_ _05621_ VPWR VGND sg13g2_nand2_1
XFILLER_14_944 VPWR VGND sg13g2_decap_8
XFILLER_40_240 VPWR VGND sg13g2_decap_8
X_10744_ _04704_ VPWR _04757_ VGND _04620_ _04636_ sg13g2_o21ai_1
X_13463_ _07111_ net1753 sipo.shift_reg\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_43_84 VPWR VGND sg13g2_decap_8
X_10675_ _04687_ VPWR _04688_ VGND fp16_res_pipe.add_renorm0.mantisa\[11\] _04644_
+ sg13g2_o21ai_1
XFILLER_9_458 VPWR VGND sg13g2_fill_1
XFILLER_13_498 VPWR VGND sg13g2_decap_4
XFILLER_127_813 VPWR VGND sg13g2_decap_8
XFILLER_126_301 VPWR VGND sg13g2_decap_8
X_13394_ VGND VPWR _07014_ net1696 _00804_ _07073_ sg13g2_a21oi_1
X_12414_ _06260_ _06258_ _06259_ VPWR VGND sg13g2_xnor2_1
X_12345_ _06191_ net1858 net1867 VPWR VGND sg13g2_nand2_1
XFILLER_126_378 VPWR VGND sg13g2_decap_4
XFILLER_126_367 VPWR VGND sg13g2_decap_8
X_12276_ _06122_ _06120_ _06121_ VPWR VGND sg13g2_nand2_1
X_14015_ VPWR _00566_ net75 VGND sg13g2_inv_1
X_11227_ net1663 _05191_ _05192_ VPWR VGND sg13g2_nor2b_2
XFILLER_4_56 VPWR VGND sg13g2_decap_8
X_11158_ _05128_ net1808 net1680 acc_sum.op_sign_logic0.mantisa_a\[9\] net1760 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_68_627 VPWR VGND sg13g2_decap_4
XFILLER_68_616 VPWR VGND sg13g2_fill_1
XFILLER_122_595 VPWR VGND sg13g2_fill_2
XFILLER_96_969 VPWR VGND sg13g2_decap_8
XFILLER_1_892 VPWR VGND sg13g2_decap_8
X_10109_ _04193_ _04192_ net1637 VPWR VGND sg13g2_nand2_1
X_11089_ _05063_ acc_sum.exp_mant_logic0.a\[9\] _05052_ net1760 acc_sum.seg_reg0.q\[24\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_64_800 VPWR VGND sg13g2_decap_8
XFILLER_48_340 VPWR VGND sg13g2_fill_1
X_14917_ _00718_ VGND VPWR _01437_ acc_sub.seg_reg0.q\[27\] clknet_leaf_51_clk sg13g2_dfrbpq_1
XFILLER_91_641 VPWR VGND sg13g2_decap_4
X_14848_ _00649_ VGND VPWR _01372_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[10\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_1
XFILLER_24_719 VPWR VGND sg13g2_fill_1
XFILLER_90_151 VPWR VGND sg13g2_decap_8
XFILLER_63_398 VPWR VGND sg13g2_fill_1
XFILLER_17_760 VPWR VGND sg13g2_fill_2
X_07320_ _01681_ _01683_ _01680_ _01480_ VPWR VGND sg13g2_nand3_1
X_14779_ _00580_ VGND VPWR _01303_ acc_sub.y\[8\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_16_292 VPWR VGND sg13g2_decap_8
XFILLER_32_741 VPWR VGND sg13g2_decap_4
XFILLER_32_752 VPWR VGND sg13g2_fill_1
X_07251_ _01620_ net1744 _01616_ _01621_ VPWR VGND sg13g2_nand3_1
X_07182_ VPWR _01554_ acc_sub.op_sign_logic0.mantisa_b\[3\] VGND sg13g2_inv_1
XFILLER_118_824 VPWR VGND sg13g2_decap_8
XFILLER_76_0 VPWR VGND sg13g2_fill_2
XFILLER_20_969 VPWR VGND sg13g2_decap_8
XFILLER_126_890 VPWR VGND sg13g2_decap_8
XFILLER_99_763 VPWR VGND sg13g2_decap_4
X_09823_ _03858_ _03855_ _03935_ VPWR VGND sg13g2_nor2_1
XFILLER_58_115 VPWR VGND sg13g2_fill_1
XFILLER_58_104 VPWR VGND sg13g2_decap_8
XFILLER_24_1009 VPWR VGND sg13g2_decap_4
XFILLER_101_757 VPWR VGND sg13g2_decap_8
XFILLER_98_284 VPWR VGND sg13g2_fill_2
XFILLER_87_958 VPWR VGND sg13g2_decap_8
XFILLER_86_457 VPWR VGND sg13g2_decap_8
X_09754_ _03870_ _03851_ _03628_ VPWR VGND sg13g2_nand2_1
XFILLER_101_768 VPWR VGND sg13g2_fill_2
XFILLER_100_267 VPWR VGND sg13g2_fill_1
XFILLER_73_107 VPWR VGND sg13g2_fill_1
XFILLER_39_362 VPWR VGND sg13g2_decap_8
X_08705_ VGND VPWR _02916_ net1817 _01336_ _02917_ sg13g2_a21oi_1
X_09685_ _03800_ _03788_ _03801_ VPWR VGND sg13g2_nor2b_1
XFILLER_67_693 VPWR VGND sg13g2_decap_8
X_08636_ _02724_ VPWR _02858_ VGND _02796_ _02793_ sg13g2_o21ai_1
Xclkbuf_leaf_93_clk clknet_5_12__leaf_clk clknet_leaf_93_clk VPWR VGND sg13g2_buf_8
XFILLER_81_151 VPWR VGND sg13g2_decap_4
XFILLER_54_387 VPWR VGND sg13g2_decap_4
XFILLER_42_538 VPWR VGND sg13g2_decap_8
XFILLER_120_56 VPWR VGND sg13g2_decap_8
X_08567_ VPWR _02791_ _02790_ VGND sg13g2_inv_1
Xfanout22 net23 net22 VPWR VGND sg13g2_buf_2
Xfanout11 net13 net11 VPWR VGND sg13g2_buf_2
X_07518_ _01839_ VPWR _01438_ VGND _01824_ net1796 sg13g2_o21ai_1
X_08498_ _02723_ VPWR _01349_ VGND _02722_ _01758_ sg13g2_o21ai_1
Xfanout33 net34 net33 VPWR VGND sg13g2_buf_2
Xfanout55 net56 net55 VPWR VGND sg13g2_buf_1
XFILLER_11_903 VPWR VGND sg13g2_decap_8
Xfanout44 net46 net44 VPWR VGND sg13g2_buf_2
X_07449_ VGND VPWR _01443_ acc_sub.reg_add_sub.q\[0\] net1895 sg13g2_or2_1
Xfanout99 net100 net99 VPWR VGND sg13g2_buf_1
Xfanout77 net80 net77 VPWR VGND sg13g2_buf_2
Xfanout88 net92 net88 VPWR VGND sg13g2_buf_2
Xfanout66 net67 net66 VPWR VGND sg13g2_buf_2
XFILLER_13_21 VPWR VGND sg13g2_decap_8
XFILLER_22_295 VPWR VGND sg13g2_decap_8
X_10460_ VPWR _04508_ _04507_ VGND sg13g2_inv_1
XFILLER_10_457 VPWR VGND sg13g2_decap_8
X_09119_ _03300_ _03299_ _03204_ VPWR VGND sg13g2_nand2b_1
XFILLER_109_835 VPWR VGND sg13g2_decap_8
XFILLER_89_14 VPWR VGND sg13g2_fill_1
XFILLER_6_439 VPWR VGND sg13g2_decap_8
XFILLER_124_816 VPWR VGND sg13g2_decap_8
X_10391_ VPWR _04441_ _04440_ VGND sg13g2_inv_1
XFILLER_123_315 VPWR VGND sg13g2_decap_8
X_12130_ _05973_ _05940_ _05976_ VPWR VGND sg13g2_nor2_1
X_12061_ VGND VPWR _05898_ _05905_ _05907_ _05906_ sg13g2_a21oi_1
XFILLER_2_645 VPWR VGND sg13g2_fill_1
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_104_584 VPWR VGND sg13g2_decap_8
X_11012_ acc_sum.op_sign_logic0.s_b acc_sum.exp_mant_logic0.b\[15\] net1813 _01103_
+ VPWR VGND sg13g2_mux2_1
XFILLER_78_936 VPWR VGND sg13g2_fill_1
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_77_468 VPWR VGND sg13g2_fill_1
XFILLER_86_980 VPWR VGND sg13g2_decap_8
X_12963_ _06733_ VPWR _06734_ VGND net1961 _06731_ sg13g2_o21ai_1
XFILLER_64_118 VPWR VGND sg13g2_decap_8
XFILLER_46_822 VPWR VGND sg13g2_decap_8
XFILLER_38_84 VPWR VGND sg13g2_decap_8
XFILLER_18_513 VPWR VGND sg13g2_decap_4
X_14702_ _00503_ VGND VPWR _01230_ acc_sum.y\[5\] clknet_leaf_39_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_84_clk clknet_5_27__leaf_clk clknet_leaf_84_clk VPWR VGND sg13g2_buf_8
XFILLER_73_663 VPWR VGND sg13g2_fill_1
X_11914_ VGND VPWR net1881 _05785_ _00996_ _05786_ sg13g2_a21oi_1
XFILLER_18_568 VPWR VGND sg13g2_fill_1
X_12894_ _06669_ _06670_ _06660_ _00901_ VPWR VGND sg13g2_nand3_1
XFILLER_45_365 VPWR VGND sg13g2_decap_8
X_14633_ _00434_ VGND VPWR _01165_ fp16_sum_pipe.add_renorm0.mantisa\[4\] clknet_leaf_108_clk
+ sg13g2_dfrbpq_2
X_11845_ VGND VPWR _05742_ _05635_ _05743_ _05636_ sg13g2_a21oi_1
X_14564_ _00365_ VGND VPWR _01100_ acc_sum.seg_reg0.q\[27\] clknet_leaf_27_clk sg13g2_dfrbpq_2
X_11776_ net1758 VPWR _05679_ VGND _05673_ _05678_ sg13g2_o21ai_1
X_14495_ _00296_ VGND VPWR _01031_ fpdiv.divider0.divisor\[6\] clknet_leaf_85_clk
+ sg13g2_dfrbpq_1
X_13515_ VPWR _00066_ net38 VGND sg13g2_inv_1
X_10727_ _04740_ net1710 VPWR VGND sg13g2_inv_2
XFILLER_70_71 VPWR VGND sg13g2_decap_4
XFILLER_127_643 VPWR VGND sg13g2_decap_8
Xclkload14 clknet_5_29__leaf_clk clkload14/Y VPWR VGND sg13g2_inv_4
Xclkload25 VPWR clkload25/Y clknet_leaf_139_clk VGND sg13g2_inv_1
XFILLER_115_816 VPWR VGND sg13g2_decap_8
Xclkload69 clknet_leaf_28_clk clkload69/Y VPWR VGND sg13g2_inv_4
Xclkload58 clkload58/Y clknet_leaf_95_clk VPWR VGND sg13g2_inv_2
X_13377_ _07065_ net1695 sipo.word\[10\] VPWR VGND sg13g2_nand2_1
Xclkload36 VPWR clkload36/Y clknet_leaf_12_clk VGND sg13g2_inv_1
Xclkload47 clknet_leaf_108_clk clkload47/X VPWR VGND sg13g2_buf_8
XFILLER_6_962 VPWR VGND sg13g2_decap_8
XFILLER_5_450 VPWR VGND sg13g2_decap_8
X_10589_ _04607_ VPWR _01142_ VGND net1934 _02260_ sg13g2_o21ai_1
XFILLER_126_175 VPWR VGND sg13g2_decap_8
XFILLER_114_326 VPWR VGND sg13g2_decap_8
X_12328_ _06174_ _06157_ _06172_ VPWR VGND sg13g2_nand2_1
X_12259_ _06094_ _06102_ _06101_ _06105_ VPWR VGND sg13g2_nand3_1
XFILLER_69_936 VPWR VGND sg13g2_decap_8
XFILLER_69_925 VPWR VGND sg13g2_fill_1
XFILLER_110_510 VPWR VGND sg13g2_decap_8
XFILLER_69_947 VPWR VGND sg13g2_fill_1
XFILLER_68_424 VPWR VGND sg13g2_decap_8
XFILLER_84_917 VPWR VGND sg13g2_decap_8
XFILLER_77_980 VPWR VGND sg13g2_fill_1
XFILLER_49_693 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_75_clk clknet_5_27__leaf_clk clknet_leaf_75_clk VPWR VGND sg13g2_buf_8
X_09470_ _03598_ acc_sub.x2\[10\] net1914 VPWR VGND sg13g2_nand2_1
XFILLER_91_482 VPWR VGND sg13g2_fill_1
XFILLER_91_471 VPWR VGND sg13g2_decap_8
XFILLER_52_836 VPWR VGND sg13g2_fill_2
XFILLER_52_825 VPWR VGND sg13g2_decap_8
XFILLER_51_313 VPWR VGND sg13g2_fill_2
XFILLER_51_346 VPWR VGND sg13g2_decap_8
X_08352_ _02595_ _02592_ _02594_ VPWR VGND sg13g2_nand2_1
X_07303_ _01669_ _01527_ _01607_ VPWR VGND sg13g2_nand2b_1
X_08283_ _02531_ net1658 fp16_sum_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
X_07234_ _01604_ VPWR _01605_ VGND _01537_ _01539_ sg13g2_o21ai_1
Xclkload8 clknet_5_17__leaf_clk clkload8/X VPWR VGND sg13g2_buf_8
XFILLER_30_1013 VPWR VGND sg13g2_fill_1
X_07165_ VPWR _01537_ acc_sub.op_sign_logic0.mantisa_a\[4\] VGND sg13g2_inv_1
XFILLER_117_175 VPWR VGND sg13g2_decap_8
XFILLER_105_304 VPWR VGND sg13g2_decap_8
XFILLER_121_819 VPWR VGND sg13g2_decap_8
XFILLER_59_28 VPWR VGND sg13g2_decap_8
XFILLER_114_860 VPWR VGND sg13g2_decap_8
XFILLER_87_744 VPWR VGND sg13g2_fill_2
XFILLER_86_210 VPWR VGND sg13g2_fill_1
XFILLER_115_56 VPWR VGND sg13g2_decap_8
X_09806_ _03920_ net1768 acc_sum.y\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_101_554 VPWR VGND sg13g2_fill_2
XFILLER_47_608 VPWR VGND sg13g2_fill_1
X_07998_ _02208_ _02264_ _02203_ _02265_ VPWR VGND _02218_ sg13g2_nand4_1
X_09737_ _03852_ VPWR _03853_ VGND _03843_ _03847_ sg13g2_o21ai_1
XFILLER_86_298 VPWR VGND sg13g2_fill_1
XFILLER_28_822 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_66_clk clknet_5_29__leaf_clk clknet_leaf_66_clk VPWR VGND sg13g2_buf_8
XFILLER_39_181 VPWR VGND sg13g2_fill_2
XFILLER_27_332 VPWR VGND sg13g2_decap_4
XFILLER_28_844 VPWR VGND sg13g2_fill_1
X_09668_ VPWR _03785_ _03783_ VGND sg13g2_inv_1
XFILLER_54_151 VPWR VGND sg13g2_decap_8
XFILLER_43_814 VPWR VGND sg13g2_decap_8
X_09599_ _03707_ _03715_ _03716_ VPWR VGND sg13g2_nor2_1
X_08619_ acc_sum.op_sign_logic0.mantisa_a\[0\] _02761_ _02841_ VPWR VGND sg13g2_nor2_2
XFILLER_42_346 VPWR VGND sg13g2_decap_4
XFILLER_27_398 VPWR VGND sg13g2_decap_8
XFILLER_70_677 VPWR VGND sg13g2_decap_8
X_11630_ _05416_ _05521_ _05535_ VPWR VGND sg13g2_nor2_1
XFILLER_24_42 VPWR VGND sg13g2_decap_8
XFILLER_11_733 VPWR VGND sg13g2_decap_4
X_13300_ acc\[3\] net1678 _07013_ VPWR VGND sg13g2_nor2_1
X_10512_ _04555_ _04443_ _04554_ VPWR VGND sg13g2_xnor2_1
X_11492_ fpdiv.divider0.divisor\[4\] fp16_res_pipe.x2\[0\] net1944 _01029_ VPWR VGND
+ sg13g2_mux2_1
X_14280_ _00081_ VGND VPWR _00831_ fp16_res_pipe.x2\[13\] clknet_leaf_16_clk sg13g2_dfrbpq_2
X_13231_ net1742 _02592_ _02580_ _06956_ VPWR VGND sg13g2_nor3_1
XFILLER_40_63 VPWR VGND sg13g2_decap_8
XFILLER_6_247 VPWR VGND sg13g2_decap_4
X_10443_ _04384_ _04491_ _04492_ VPWR VGND sg13g2_nor2_1
XFILLER_124_613 VPWR VGND sg13g2_fill_2
XFILLER_109_687 VPWR VGND sg13g2_decap_8
XFILLER_108_153 VPWR VGND sg13g2_decap_8
X_10374_ VPWR _04424_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[3\] VGND sg13g2_inv_1
XFILLER_3_910 VPWR VGND sg13g2_decap_8
XFILLER_124_646 VPWR VGND sg13g2_decap_8
XFILLER_123_112 VPWR VGND sg13g2_decap_8
XFILLER_97_508 VPWR VGND sg13g2_fill_1
X_12113_ _05959_ net1857 net1865 VPWR VGND sg13g2_nand2_1
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_124_679 VPWR VGND sg13g2_decap_8
XFILLER_111_307 VPWR VGND sg13g2_fill_2
XFILLER_105_882 VPWR VGND sg13g2_fill_1
X_13093_ VGND VPWR _06802_ _06765_ _06854_ _06835_ sg13g2_a21oi_1
XFILLER_3_987 VPWR VGND sg13g2_decap_8
XFILLER_123_189 VPWR VGND sg13g2_decap_8
XFILLER_120_841 VPWR VGND sg13g2_decap_8
X_12044_ _05890_ net1859 net1863 VPWR VGND sg13g2_nand2_1
XFILLER_2_486 VPWR VGND sg13g2_decap_8
XFILLER_78_788 VPWR VGND sg13g2_fill_2
XFILLER_38_619 VPWR VGND sg13g2_fill_2
XFILLER_93_736 VPWR VGND sg13g2_decap_8
XFILLER_65_427 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_57_clk clknet_5_25__leaf_clk clknet_leaf_57_clk VPWR VGND sg13g2_buf_8
X_13995_ VPWR _00546_ net15 VGND sg13g2_inv_1
X_12946_ _06718_ net1910 fp16_res_pipe.y\[2\] VPWR VGND sg13g2_nand2_2
XFILLER_45_140 VPWR VGND sg13g2_decap_8
X_12877_ VPWR _06655_ fpmul.reg_p_out\[8\] VGND sg13g2_inv_1
X_14616_ _00417_ VGND VPWR _01148_ fp16_sum_pipe.exp_mant_logic0.a\[11\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_2
X_11828_ net1837 _05727_ _05722_ _05728_ VPWR VGND sg13g2_nand3_1
X_14547_ _00348_ VGND VPWR _01083_ acc_sum.op_sign_logic0.mantisa_b\[10\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_81_70 VPWR VGND sg13g2_decap_8
XFILLER_14_571 VPWR VGND sg13g2_fill_1
XFILLER_41_390 VPWR VGND sg13g2_decap_8
X_11759_ net1838 fp16_sum_pipe.add_renorm0.exp\[0\] _05663_ VPWR VGND sg13g2_nor2_1
XFILLER_119_429 VPWR VGND sg13g2_fill_2
Xclkload103 clknet_leaf_77_clk clkload103/Y VPWR VGND sg13g2_inv_4
X_14478_ _00279_ VGND VPWR _01016_ add_result\[3\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_127_451 VPWR VGND sg13g2_decap_8
XFILLER_127_440 VPWR VGND sg13g2_fill_1
Xclkload114 clkload114/Y clknet_leaf_73_clk VPWR VGND sg13g2_inv_2
X_13429_ _07093_ VPWR _00789_ VGND _07010_ net1719 sg13g2_o21ai_1
Xplace1904 net1903 net1904 VPWR VGND sg13g2_buf_1
Xplace1915 net1913 net1915 VPWR VGND sg13g2_buf_2
Xplace1926 net1925 net1926 VPWR VGND sg13g2_buf_2
XFILLER_114_112 VPWR VGND sg13g2_decap_8
Xplace1948 net1944 net1948 VPWR VGND sg13g2_buf_2
Xplace1937 fpdiv.reg1en.d\[0\] net1937 VPWR VGND sg13g2_buf_1
Xplace1959 net1958 net1959 VPWR VGND sg13g2_buf_1
XFILLER_115_679 VPWR VGND sg13g2_decap_8
X_08970_ acc_sub.add_renorm0.exp\[3\] net1699 _03156_ VPWR VGND sg13g2_nor2_1
XFILLER_69_733 VPWR VGND sg13g2_fill_1
XFILLER_68_210 VPWR VGND sg13g2_decap_8
XFILLER_39_0 VPWR VGND sg13g2_decap_8
X_07921_ _02193_ _02195_ _02196_ VPWR VGND sg13g2_nor2_1
XFILLER_111_852 VPWR VGND sg13g2_decap_8
X_07852_ _02145_ _02146_ _02147_ VPWR VGND _02140_ sg13g2_nand3b_1
XFILLER_96_541 VPWR VGND sg13g2_fill_1
XFILLER_57_917 VPWR VGND sg13g2_decap_4
Xinput1 mosi net1 VPWR VGND sg13g2_buf_2
XFILLER_84_736 VPWR VGND sg13g2_decap_8
XFILLER_69_799 VPWR VGND sg13g2_decap_4
X_09522_ _03638_ VPWR _03639_ VGND _03634_ _03637_ sg13g2_o21ai_1
X_07783_ _02083_ acc_sub.exp_mant_logic0.b\[4\] net1651 net1685 acc_sub.exp_mant_logic0.b\[3\]
+ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_48_clk clknet_5_20__leaf_clk clknet_leaf_48_clk VPWR VGND sg13g2_buf_8
XFILLER_84_758 VPWR VGND sg13g2_decap_8
XFILLER_71_408 VPWR VGND sg13g2_fill_2
XFILLER_52_611 VPWR VGND sg13g2_fill_2
XFILLER_91_290 VPWR VGND sg13g2_decap_4
XFILLER_80_953 VPWR VGND sg13g2_decap_4
XFILLER_36_184 VPWR VGND sg13g2_decap_8
X_09453_ _03587_ VPWR _01258_ VGND net1832 _03586_ sg13g2_o21ai_1
X_08404_ _02566_ _02637_ _02639_ _02640_ VPWR VGND sg13g2_nor3_1
X_09384_ _03532_ net1770 fp16_res_pipe.add_renorm0.mantisa\[6\] VPWR VGND sg13g2_nand2_1
X_08335_ VPWR _02580_ _02579_ VGND sg13g2_inv_1
XFILLER_61_18 VPWR VGND sg13g2_decap_4
X_08266_ _02516_ fp16_sum_pipe.exp_mant_logic0.b\[1\] _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[4\]
+ net1778 VPWR VGND sg13g2_a22oi_1
X_07217_ _01543_ _01566_ _01581_ _01589_ VPWR VGND _01588_ sg13g2_nand4_1
XFILLER_117_7 VPWR VGND sg13g2_decap_8
X_08197_ _02454_ _02448_ _02453_ VPWR VGND sg13g2_nand2_1
XFILLER_119_996 VPWR VGND sg13g2_decap_8
X_07148_ acc_sub.op_sign_logic0.mantisa_a\[7\] _01519_ _01520_ VPWR VGND sg13g2_nor2_1
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_3_217 VPWR VGND sg13g2_fill_2
XFILLER_121_616 VPWR VGND sg13g2_fill_1
XFILLER_105_156 VPWR VGND sg13g2_decap_8
XFILLER_105_145 VPWR VGND sg13g2_fill_2
XFILLER_10_77 VPWR VGND sg13g2_decap_8
XFILLER_126_77 VPWR VGND sg13g2_decap_8
XFILLER_121_649 VPWR VGND sg13g2_decap_8
XFILLER_120_126 VPWR VGND sg13g2_decap_8
XFILLER_86_26 VPWR VGND sg13g2_decap_8
X_10090_ _04175_ net1662 _04146_ VPWR VGND sg13g2_nand2_2
XFILLER_87_541 VPWR VGND sg13g2_decap_8
XFILLER_75_703 VPWR VGND sg13g2_decap_8
XFILLER_0_968 VPWR VGND sg13g2_decap_8
XFILLER_102_885 VPWR VGND sg13g2_decap_4
XFILLER_101_373 VPWR VGND sg13g2_fill_1
XFILLER_59_276 VPWR VGND sg13g2_decap_8
XFILLER_47_416 VPWR VGND sg13g2_decap_8
XFILLER_19_42 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_39_clk clknet_5_21__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_74_257 VPWR VGND sg13g2_decap_8
X_12800_ _06583_ _06582_ net1923 _06584_ VPWR VGND sg13g2_a21o_1
X_13780_ VPWR _00331_ net124 VGND sg13g2_inv_1
XFILLER_56_983 VPWR VGND sg13g2_decap_8
XFILLER_27_140 VPWR VGND sg13g2_decap_4
X_10992_ _04982_ fp16_res_pipe.x2\[8\] net1932 VPWR VGND sg13g2_nand2_1
X_12731_ _06513_ VPWR _06535_ VGND net1734 _06534_ sg13g2_o21ai_1
XFILLER_55_493 VPWR VGND sg13g2_decap_8
XFILLER_55_482 VPWR VGND sg13g2_decap_8
XFILLER_16_847 VPWR VGND sg13g2_decap_8
X_12662_ _06478_ _06366_ VPWR VGND sg13g2_inv_2
XFILLER_71_986 VPWR VGND sg13g2_decap_4
XFILLER_43_666 VPWR VGND sg13g2_fill_2
XFILLER_37_1008 VPWR VGND sg13g2_decap_4
XFILLER_35_63 VPWR VGND sg13g2_decap_8
X_14401_ _00202_ VGND VPWR _00940_ div_result\[14\] clknet_leaf_89_clk sg13g2_dfrbpq_1
XFILLER_70_474 VPWR VGND sg13g2_decap_4
X_11613_ net1840 fp16_sum_pipe.add_renorm0.mantisa\[0\] _05518_ VPWR VGND sg13g2_nor2_1
X_12593_ fpdiv.reg_b_out\[12\] _05361_ _06409_ VPWR VGND sg13g2_nor2_1
XFILLER_11_530 VPWR VGND sg13g2_decap_8
X_14332_ _00133_ VGND VPWR _00874_ piso.tx_bit_counter\[1\] clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_11_552 VPWR VGND sg13g2_fill_1
X_11544_ VPWR _05449_ _05448_ VGND sg13g2_inv_1
XFILLER_125_900 VPWR VGND sg13g2_decap_8
XFILLER_100_1000 VPWR VGND sg13g2_decap_8
X_11475_ VPWR _05389_ fpdiv.reg_b_out\[8\] VGND sg13g2_inv_1
X_14263_ _00064_ VGND VPWR _00814_ acc_sub.x2\[12\] clknet_leaf_127_clk sg13g2_dfrbpq_2
XFILLER_51_95 VPWR VGND sg13g2_decap_8
XFILLER_124_410 VPWR VGND sg13g2_fill_1
X_13214_ _06943_ sipo.bit_counter\[4\] _00854_ VPWR VGND sg13g2_nor2b_1
XFILLER_7_578 VPWR VGND sg13g2_fill_2
X_10426_ _04475_ _04474_ _04473_ VPWR VGND sg13g2_nand2b_1
X_14194_ VPWR _00745_ net91 VGND sg13g2_inv_1
XFILLER_125_977 VPWR VGND sg13g2_decap_8
X_13145_ VGND VPWR _06891_ _06882_ _06894_ piso.tx_bit_counter\[0\] sg13g2_a21oi_1
X_10357_ _04407_ _04406_ VPWR VGND sg13g2_inv_2
XFILLER_97_349 VPWR VGND sg13g2_fill_1
X_13076_ _06842_ VPWR _00891_ VGND net1861 _06599_ sg13g2_o21ai_1
XFILLER_2_272 VPWR VGND sg13g2_decap_8
X_10288_ _04351_ _04356_ _04357_ VPWR VGND _04350_ sg13g2_nand3b_1
XFILLER_32_7 VPWR VGND sg13g2_decap_8
XFILLER_111_159 VPWR VGND sg13g2_decap_8
XFILLER_78_563 VPWR VGND sg13g2_fill_1
X_12027_ net1873 _05874_ _05875_ VPWR VGND _05843_ sg13g2_nand3b_1
XFILLER_93_522 VPWR VGND sg13g2_decap_4
XFILLER_78_585 VPWR VGND sg13g2_fill_2
XFILLER_93_566 VPWR VGND sg13g2_decap_8
XFILLER_53_419 VPWR VGND sg13g2_fill_2
X_13978_ VPWR _00529_ net26 VGND sg13g2_inv_1
XFILLER_19_685 VPWR VGND sg13g2_decap_8
X_12929_ _06703_ net1717 _00009_ VPWR VGND sg13g2_nand2_1
XFILLER_74_780 VPWR VGND sg13g2_decap_4
XFILLER_62_975 VPWR VGND sg13g2_decap_8
XFILLER_34_666 VPWR VGND sg13g2_decap_8
XFILLER_33_154 VPWR VGND sg13g2_fill_2
XFILLER_21_316 VPWR VGND sg13g2_decap_4
XFILLER_33_198 VPWR VGND sg13g2_decap_8
XFILLER_119_259 VPWR VGND sg13g2_decap_8
X_08051_ _02316_ VPWR _02317_ VGND _02217_ net1692 sg13g2_o21ai_1
XFILLER_116_933 VPWR VGND sg13g2_decap_8
Xplace1701 _06567_ net1701 VPWR VGND sg13g2_buf_2
XFILLER_115_421 VPWR VGND sg13g2_fill_2
Xplace1734 _06366_ net1734 VPWR VGND sg13g2_buf_2
Xplace1723 _07027_ net1723 VPWR VGND sg13g2_buf_2
Xplace1712 _06907_ net1712 VPWR VGND sg13g2_buf_2
Xplace1745 _04268_ net1745 VPWR VGND sg13g2_buf_2
Xplace1767 _03983_ net1767 VPWR VGND sg13g2_buf_2
Xplace1756 _05573_ net1756 VPWR VGND sg13g2_buf_2
Xplace1778 net1777 net1778 VPWR VGND sg13g2_buf_1
Xplace1789 net1788 net1789 VPWR VGND sg13g2_buf_2
X_08953_ acc_sub.add_renorm0.exp\[1\] acc_sub.add_renorm0.exp\[0\] acc_sub.add_renorm0.exp\[2\]
+ _03139_ VPWR VGND sg13g2_nand3_1
XFILLER_88_349 VPWR VGND sg13g2_fill_2
X_07904_ _02179_ fp16_sum_pipe.reg1en.q\[0\] VPWR VGND sg13g2_inv_2
X_08884_ VGND VPWR _03059_ _03027_ _03071_ _03070_ sg13g2_a21oi_1
XFILLER_69_574 VPWR VGND sg13g2_decap_8
XFILLER_29_416 VPWR VGND sg13g2_fill_1
XFILLER_29_427 VPWR VGND sg13g2_fill_2
XFILLER_110_181 VPWR VGND sg13g2_fill_2
X_07835_ _02131_ _01949_ acc_sub.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
X_07766_ _02068_ net1651 net1794 VPWR VGND sg13g2_nand2_1
XFILLER_112_35 VPWR VGND sg13g2_decap_8
X_09505_ VPWR _03622_ _03621_ VGND sg13g2_inv_1
XFILLER_38_994 VPWR VGND sg13g2_decap_8
X_07697_ _02005_ _01940_ _01928_ VPWR VGND sg13g2_nand2_1
X_09436_ _03576_ fp16_res_pipe.add_renorm0.exp\[6\] VPWR VGND sg13g2_inv_2
XFILLER_25_655 VPWR VGND sg13g2_decap_8
XFILLER_80_783 VPWR VGND sg13g2_decap_4
XFILLER_12_316 VPWR VGND sg13g2_decap_4
XFILLER_8_309 VPWR VGND sg13g2_fill_2
X_09367_ _03517_ _03475_ fp16_res_pipe.reg2en.q\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_24_198 VPWR VGND sg13g2_fill_1
X_08318_ _02560_ _02562_ _02563_ VPWR VGND sg13g2_nor2_2
X_09298_ _03451_ _03438_ _03442_ _03452_ VPWR VGND _03390_ sg13g2_nand4_1
X_08249_ _02497_ _02498_ _02499_ _02500_ VPWR VGND sg13g2_nor3_1
XFILLER_20_371 VPWR VGND sg13g2_decap_8
XFILLER_21_21 VPWR VGND sg13g2_decap_8
XFILLER_107_922 VPWR VGND sg13g2_decap_8
XFILLER_4_504 VPWR VGND sg13g2_decap_8
XFILLER_119_793 VPWR VGND sg13g2_decap_8
X_11260_ _05223_ net1655 acc_sum.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_122_903 VPWR VGND sg13g2_decap_8
XFILLER_107_999 VPWR VGND sg13g2_decap_8
XFILLER_106_476 VPWR VGND sg13g2_decap_8
X_11191_ _01092_ _05158_ _05159_ VPWR VGND sg13g2_nand2_1
X_10211_ _04286_ _04285_ net1636 VPWR VGND sg13g2_nand2_1
XFILLER_121_435 VPWR VGND sg13g2_decap_4
XFILLER_79_327 VPWR VGND sg13g2_fill_2
XFILLER_0_721 VPWR VGND sg13g2_decap_8
X_14950_ _00751_ VGND VPWR _01470_ acc_sub.add_renorm0.exp\[2\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
XFILLER_94_308 VPWR VGND sg13g2_decap_8
XFILLER_0_743 VPWR VGND sg13g2_decap_8
X_10073_ _04160_ net1688 net1828 VPWR VGND sg13g2_nand2_1
X_14881_ _00682_ VGND VPWR _01401_ acc_sub.exp_mant_logic0.b\[7\] clknet_leaf_61_clk
+ sg13g2_dfrbpq_1
XFILLER_47_235 VPWR VGND sg13g2_fill_2
X_13901_ VPWR _00452_ net11 VGND sg13g2_inv_1
XFILLER_75_577 VPWR VGND sg13g2_decap_4
XFILLER_47_268 VPWR VGND sg13g2_fill_1
X_13832_ VPWR _00383_ net52 VGND sg13g2_inv_1
XFILLER_28_460 VPWR VGND sg13g2_fill_2
XFILLER_29_983 VPWR VGND sg13g2_decap_8
X_13763_ VPWR _00314_ net117 VGND sg13g2_inv_1
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_44_942 VPWR VGND sg13g2_decap_8
XFILLER_28_482 VPWR VGND sg13g2_decap_8
X_12714_ VPWR _06520_ div_result\[4\] VGND sg13g2_inv_1
X_10975_ VGND VPWR _04973_ net1835 _01123_ _04974_ sg13g2_a21oi_1
XFILLER_44_953 VPWR VGND sg13g2_fill_2
XFILLER_15_121 VPWR VGND sg13g2_fill_1
XFILLER_71_794 VPWR VGND sg13g2_fill_1
X_13694_ VPWR _00245_ net66 VGND sg13g2_inv_1
XFILLER_15_154 VPWR VGND sg13g2_decap_8
XFILLER_16_688 VPWR VGND sg13g2_fill_1
XFILLER_16_699 VPWR VGND sg13g2_decap_8
Xclkbuf_5_0__f_clk clknet_4_0_0_clk clknet_5_0__leaf_clk VPWR VGND sg13g2_buf_8
X_12645_ _06420_ _06460_ _06461_ VPWR VGND sg13g2_nor2_1
XFILLER_62_61 VPWR VGND sg13g2_fill_1
XFILLER_31_658 VPWR VGND sg13g2_fill_2
X_12576_ _06391_ _06390_ _06392_ VPWR VGND sg13g2_xor2_1
XFILLER_62_94 VPWR VGND sg13g2_decap_4
XFILLER_50_1005 VPWR VGND sg13g2_decap_8
XFILLER_8_832 VPWR VGND sg13g2_decap_8
XFILLER_12_883 VPWR VGND sg13g2_decap_8
XFILLER_30_179 VPWR VGND sg13g2_fill_2
X_14315_ _00116_ VGND VPWR _00858_ sipo.word\[3\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_11_382 VPWR VGND sg13g2_fill_2
X_11527_ VPWR _05432_ fp16_sum_pipe.add_renorm0.mantisa\[3\] VGND sg13g2_inv_1
XFILLER_7_375 VPWR VGND sg13g2_fill_1
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_116_229 VPWR VGND sg13g2_decap_8
X_11458_ _05381_ VPWR _01047_ VGND net1947 _05380_ sg13g2_o21ai_1
X_14246_ _00047_ VGND VPWR _00797_ instr\[11\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_125_774 VPWR VGND sg13g2_decap_8
XFILLER_113_914 VPWR VGND sg13g2_decap_8
X_11389_ _05338_ net1707 fpdiv.div_out\[11\] VPWR VGND sg13g2_nand2_1
X_14177_ VPWR _00728_ net127 VGND sg13g2_inv_1
X_10409_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[10\] _02259_ _04459_ VPWR VGND sg13g2_nor2_1
XFILLER_124_273 VPWR VGND sg13g2_decap_8
X_13128_ _06880_ VPWR _06881_ VGND _06564_ _06558_ sg13g2_o21ai_1
XFILLER_97_135 VPWR VGND sg13g2_fill_2
XFILLER_121_980 VPWR VGND sg13g2_decap_8
XFILLER_112_479 VPWR VGND sg13g2_decap_8
XFILLER_94_820 VPWR VGND sg13g2_fill_1
X_13059_ fpmul.seg_reg0.q\[50\] _06824_ _06826_ _06827_ VPWR VGND sg13g2_nor3_1
XFILLER_39_747 VPWR VGND sg13g2_decap_8
X_07620_ _01819_ _01933_ _01934_ VPWR VGND sg13g2_nor2_1
XFILLER_19_460 VPWR VGND sg13g2_fill_2
XFILLER_26_419 VPWR VGND sg13g2_decap_8
X_07551_ _01727_ _01729_ _01725_ _01866_ VPWR VGND _01731_ sg13g2_nand4_1
XFILLER_81_569 VPWR VGND sg13g2_decap_4
XFILLER_62_761 VPWR VGND sg13g2_decap_4
XFILLER_50_901 VPWR VGND sg13g2_fill_2
XFILLER_35_953 VPWR VGND sg13g2_decap_8
XFILLER_107_1006 VPWR VGND sg13g2_decap_8
X_07482_ acc_sub.exp_mant_logic0.a\[10\] _01804_ _01805_ VPWR VGND sg13g2_nor2_1
X_09221_ _03375_ _03372_ fp16_res_pipe.op_sign_logic0.mantisa_b\[9\] VPWR VGND sg13g2_nand2_1
X_09152_ _03325_ net1773 acc_sub.y\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_21_168 VPWR VGND sg13g2_fill_2
X_08103_ _02367_ net1639 _02366_ VPWR VGND sg13g2_nand2_1
X_09083_ _03267_ _03209_ _03183_ VPWR VGND sg13g2_nand2_1
XFILLER_108_719 VPWR VGND sg13g2_fill_1
X_08034_ _02299_ _02201_ _02300_ VPWR VGND sg13g2_xor2_1
XFILLER_115_284 VPWR VGND sg13g2_fill_2
XFILLER_115_273 VPWR VGND sg13g2_decap_8
XFILLER_107_35 VPWR VGND sg13g2_decap_8
XFILLER_104_936 VPWR VGND sg13g2_decap_8
XFILLER_89_636 VPWR VGND sg13g2_fill_2
XFILLER_115_295 VPWR VGND sg13g2_fill_2
XFILLER_103_457 VPWR VGND sg13g2_decap_8
XFILLER_89_669 VPWR VGND sg13g2_fill_2
XFILLER_67_39 VPWR VGND sg13g2_decap_4
XFILLER_67_28 VPWR VGND sg13g2_fill_2
X_08936_ _03060_ _03023_ _03123_ VPWR VGND sg13g2_nor2b_1
XFILLER_88_179 VPWR VGND sg13g2_decap_4
XFILLER_85_820 VPWR VGND sg13g2_fill_2
X_08867_ _03048_ _03053_ _03054_ VPWR VGND sg13g2_nor2_2
XFILLER_69_393 VPWR VGND sg13g2_decap_8
XFILLER_123_56 VPWR VGND sg13g2_decap_8
X_07818_ _02115_ net1649 acc_sub.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_84_352 VPWR VGND sg13g2_decap_8
XFILLER_57_566 VPWR VGND sg13g2_decap_8
XFILLER_57_555 VPWR VGND sg13g2_fill_1
X_08798_ VPWR _02985_ acc_sub.add_renorm0.mantisa\[2\] VGND sg13g2_inv_1
XFILLER_84_396 VPWR VGND sg13g2_decap_8
XFILLER_83_38 VPWR VGND sg13g2_decap_8
XFILLER_45_739 VPWR VGND sg13g2_fill_2
X_07749_ _02053_ VPWR _01421_ VGND net1796 _02042_ sg13g2_o21ai_1
XFILLER_72_558 VPWR VGND sg13g2_decap_4
XFILLER_37_290 VPWR VGND sg13g2_decap_8
XFILLER_16_21 VPWR VGND sg13g2_decap_8
XFILLER_26_975 VPWR VGND sg13g2_decap_8
X_10760_ _04773_ _04772_ fp16_res_pipe.y\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_13_614 VPWR VGND sg13g2_decap_8
X_09419_ _03462_ net1738 _03563_ VPWR VGND sg13g2_and2_1
XFILLER_12_135 VPWR VGND sg13g2_fill_2
XFILLER_13_658 VPWR VGND sg13g2_decap_8
X_10691_ VPWR _04704_ _04632_ VGND sg13g2_inv_1
X_12430_ _06260_ _06261_ _06276_ VPWR VGND sg13g2_nor2_1
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_21_680 VPWR VGND sg13g2_fill_2
XFILLER_32_42 VPWR VGND sg13g2_decap_8
X_12361_ VGND VPWR _06202_ _06204_ _06207_ _06206_ sg13g2_a21oi_1
X_14100_ VPWR _00651_ net42 VGND sg13g2_inv_1
X_12292_ _06138_ _06137_ _05974_ VPWR VGND sg13g2_nand2_1
X_11312_ _05269_ net1634 _05268_ VPWR VGND sg13g2_nand2_1
XFILLER_5_857 VPWR VGND sg13g2_decap_8
X_14031_ VPWR _00582_ net106 VGND sg13g2_inv_1
XFILLER_107_752 VPWR VGND sg13g2_decap_8
XFILLER_106_0 VPWR VGND sg13g2_decap_8
X_11243_ _05204_ _05206_ _05207_ VPWR VGND sg13g2_nor2_1
XFILLER_121_210 VPWR VGND sg13g2_decap_8
XFILLER_110_906 VPWR VGND sg13g2_decap_8
XFILLER_79_135 VPWR VGND sg13g2_decap_8
X_11174_ _05143_ _05141_ VPWR VGND sg13g2_inv_2
XFILLER_0_540 VPWR VGND sg13g2_decap_8
XFILLER_122_777 VPWR VGND sg13g2_decap_8
XFILLER_94_105 VPWR VGND sg13g2_decap_4
XFILLER_88_680 VPWR VGND sg13g2_decap_8
XFILLER_0_551 VPWR VGND sg13g2_fill_2
X_10125_ _01206_ _04206_ _04207_ VPWR VGND sg13g2_nand2_1
X_14933_ _00734_ VGND VPWR _01453_ acc_sub.exp_mant_logic0.a\[1\] clknet_5_28__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_48_544 VPWR VGND sg13g2_decap_8
XFILLER_0_584 VPWR VGND sg13g2_decap_8
X_10056_ _04143_ _04122_ _04144_ VPWR VGND sg13g2_nor2_1
XFILLER_48_566 VPWR VGND sg13g2_fill_2
XFILLER_75_374 VPWR VGND sg13g2_decap_8
X_14864_ _00665_ VGND VPWR _01388_ fp16_sum_pipe.seg_reg0.q\[26\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_1
X_13815_ VPWR _00366_ net77 VGND sg13g2_inv_1
X_14795_ _00596_ VGND VPWR _01319_ acc_sum.exp_mant_logic0.a\[8\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
XFILLER_17_975 VPWR VGND sg13g2_decap_8
XFILLER_32_901 VPWR VGND sg13g2_decap_8
XFILLER_90_388 VPWR VGND sg13g2_decap_8
X_13746_ VPWR _00297_ net123 VGND sg13g2_inv_1
XFILLER_16_474 VPWR VGND sg13g2_decap_8
XFILLER_16_485 VPWR VGND sg13g2_fill_2
X_10958_ VGND VPWR _04748_ _04865_ _04963_ fp16_res_pipe.seg_reg1.q\[21\] sg13g2_a21oi_1
XFILLER_71_580 VPWR VGND sg13g2_decap_8
X_13677_ VPWR _00228_ net122 VGND sg13g2_inv_1
XFILLER_43_282 VPWR VGND sg13g2_decap_8
X_12628_ _06444_ net1852 fpdiv.div_out\[6\] VPWR VGND sg13g2_nand2_1
X_10889_ _04897_ _04899_ _04896_ _04900_ VPWR VGND sg13g2_nand3_1
XFILLER_32_978 VPWR VGND sg13g2_decap_8
X_12559_ _06374_ _06373_ _06375_ VPWR VGND sg13g2_xor2_1
XFILLER_8_684 VPWR VGND sg13g2_decap_8
XFILLER_7_172 VPWR VGND sg13g2_fill_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
X_14229_ _00030_ VGND VPWR _00780_ sipo.shift_reg\[10\] clknet_leaf_10_clk sg13g2_dfrbpq_1
XFILLER_7_194 VPWR VGND sg13g2_decap_4
XFILLER_112_243 VPWR VGND sg13g2_decap_8
XFILLER_101_906 VPWR VGND sg13g2_decap_8
XFILLER_113_788 VPWR VGND sg13g2_decap_8
XFILLER_112_254 VPWR VGND sg13g2_fill_2
X_09770_ net1769 _03876_ _03885_ _03886_ VPWR VGND sg13g2_nor3_1
XFILLER_98_488 VPWR VGND sg13g2_fill_2
XFILLER_21_0 VPWR VGND sg13g2_decap_8
X_08721_ _02927_ VPWR _01330_ VGND net1815 _02926_ sg13g2_o21ai_1
XFILLER_67_831 VPWR VGND sg13g2_fill_2
XFILLER_94_672 VPWR VGND sg13g2_fill_1
X_08652_ _02872_ _02865_ _02787_ VPWR VGND sg13g2_nand2_1
XFILLER_82_812 VPWR VGND sg13g2_fill_1
XFILLER_67_875 VPWR VGND sg13g2_fill_2
XFILLER_66_363 VPWR VGND sg13g2_fill_1
X_07603_ VGND VPWR net1686 _01915_ _01917_ _01916_ sg13g2_a21oi_1
XFILLER_82_834 VPWR VGND sg13g2_fill_2
XFILLER_39_588 VPWR VGND sg13g2_decap_8
X_08583_ acc_sum.add_renorm0.mantisa\[11\] _02806_ VPWR VGND sg13g2_inv_4
XFILLER_93_193 VPWR VGND sg13g2_decap_8
XFILLER_82_856 VPWR VGND sg13g2_fill_2
X_07534_ _01854_ net1782 acc_sub.seg_reg0.q\[26\] VPWR VGND sg13g2_nand2_1
XFILLER_23_912 VPWR VGND sg13g2_decap_8
X_07465_ acc_sub.exp_mant_logic0.b\[14\] _01725_ _01788_ VPWR VGND sg13g2_nor2_1
X_09204_ VPWR _03359_ fp16_res_pipe.seg_reg1.q\[21\] VGND sg13g2_inv_1
XFILLER_23_989 VPWR VGND sg13g2_decap_8
X_07396_ _01739_ acc_sub.exp_mant_logic0.a\[7\] VPWR VGND sg13g2_inv_2
XFILLER_108_516 VPWR VGND sg13g2_fill_1
X_09135_ _03314_ VPWR _01303_ VGND net1801 _03305_ sg13g2_o21ai_1
X_09066_ VPWR _03251_ _03210_ VGND sg13g2_inv_1
XFILLER_123_508 VPWR VGND sg13g2_fill_2
XFILLER_118_56 VPWR VGND sg13g2_decap_8
X_08017_ VPWR _02283_ _02282_ VGND sg13g2_inv_1
XFILLER_104_722 VPWR VGND sg13g2_decap_8
XFILLER_78_38 VPWR VGND sg13g2_decap_8
XFILLER_78_16 VPWR VGND sg13g2_decap_8
XFILLER_2_849 VPWR VGND sg13g2_decap_8
XFILLER_103_232 VPWR VGND sg13g2_decap_8
XFILLER_103_210 VPWR VGND sg13g2_decap_4
XFILLER_1_359 VPWR VGND sg13g2_decap_8
XFILLER_104_799 VPWR VGND sg13g2_decap_4
XFILLER_103_254 VPWR VGND sg13g2_fill_1
X_09968_ _04061_ fp16_res_pipe.exp_mant_logic0.a\[10\] _04056_ net1765 fp16_res_pipe.seg_reg0.q\[25\]
+ VPWR VGND sg13g2_a22oi_1
X_08919_ _03013_ VPWR _03106_ VGND _02994_ _03009_ sg13g2_o21ai_1
XFILLER_100_972 VPWR VGND sg13g2_decap_8
XFILLER_94_37 VPWR VGND sg13g2_fill_1
XFILLER_92_609 VPWR VGND sg13g2_decap_8
XFILLER_73_812 VPWR VGND sg13g2_decap_8
X_11930_ VPWR _05797_ fpmul.seg_reg0.q\[36\] VGND sg13g2_inv_1
X_09899_ fp16_res_pipe.exp_mant_logic0.a\[12\] _03995_ _03996_ VPWR VGND sg13g2_nor2_2
XFILLER_85_694 VPWR VGND sg13g2_decap_8
XFILLER_57_396 VPWR VGND sg13g2_fill_2
XFILLER_17_227 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_17_238 VPWR VGND sg13g2_fill_2
X_11861_ VGND VPWR _05757_ _05636_ _05758_ net1758 sg13g2_a21oi_1
XFILLER_72_366 VPWR VGND sg13g2_decap_8
X_13600_ VPWR _00151_ net59 VGND sg13g2_inv_1
XFILLER_60_528 VPWR VGND sg13g2_decap_8
X_11792_ _05648_ _05693_ _05694_ VPWR VGND _05692_ sg13g2_nand3b_1
X_14580_ _00381_ VGND VPWR _01112_ fp16_sum_pipe.exp_mant_logic0.b\[7\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_1
XFILLER_14_923 VPWR VGND sg13g2_decap_8
X_10812_ _04824_ fp16_res_pipe.add_renorm0.exp\[1\] _04823_ VPWR VGND sg13g2_xnor2_1
X_13531_ VPWR _00082_ net37 VGND sg13g2_inv_1
X_10743_ _04756_ _04626_ _04705_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_63 VPWR VGND sg13g2_decap_8
XFILLER_13_477 VPWR VGND sg13g2_decap_8
X_13462_ _07110_ VPWR _00773_ VGND _06935_ net1753 sg13g2_o21ai_1
XFILLER_40_263 VPWR VGND sg13g2_decap_8
X_10674_ _04687_ fp16_res_pipe.add_renorm0.mantisa\[11\] fp16_res_pipe.add_renorm0.mantisa\[8\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_9_437 VPWR VGND sg13g2_fill_2
XFILLER_9_448 VPWR VGND sg13g2_fill_1
X_13393_ acc_sub.x2\[2\] net1696 _07073_ VPWR VGND sg13g2_nor2_1
X_12413_ _06042_ _06037_ _06259_ VPWR VGND sg13g2_and2_1
X_12344_ VPWR _06190_ _06189_ VGND sg13g2_inv_1
XFILLER_5_621 VPWR VGND sg13g2_fill_2
XFILLER_127_869 VPWR VGND sg13g2_decap_8
X_14014_ VPWR _00565_ net75 VGND sg13g2_inv_1
X_12275_ VPWR _06121_ _05971_ VGND sg13g2_inv_1
XFILLER_4_175 VPWR VGND sg13g2_decap_8
XFILLER_107_593 VPWR VGND sg13g2_decap_8
X_11226_ _05134_ _05144_ _05191_ VPWR VGND sg13g2_nor2_1
XFILLER_4_35 VPWR VGND sg13g2_decap_8
XFILLER_110_725 VPWR VGND sg13g2_decap_8
XFILLER_96_948 VPWR VGND sg13g2_decap_8
XFILLER_68_60 VPWR VGND sg13g2_decap_8
X_11157_ _05127_ _05046_ _05126_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_871 VPWR VGND sg13g2_decap_8
X_10108_ _04187_ _04191_ _04185_ _04192_ VPWR VGND sg13g2_nand3_1
X_11088_ _05061_ _05062_ _05060_ _01098_ VPWR VGND sg13g2_nand3_1
X_14916_ _00717_ VGND VPWR _01436_ acc_sub.seg_reg0.q\[26\] clknet_leaf_50_clk sg13g2_dfrbpq_1
XFILLER_48_385 VPWR VGND sg13g2_decap_4
X_10039_ _04127_ net1746 _04126_ net1688 net1827 VPWR VGND sg13g2_a22oi_1
XFILLER_91_664 VPWR VGND sg13g2_fill_1
XFILLER_91_653 VPWR VGND sg13g2_decap_8
XFILLER_90_141 VPWR VGND sg13g2_fill_2
XFILLER_90_130 VPWR VGND sg13g2_decap_4
XFILLER_84_81 VPWR VGND sg13g2_decap_4
X_14847_ _00648_ VGND VPWR _01371_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[9\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
XFILLER_24_709 VPWR VGND sg13g2_decap_4
XFILLER_63_377 VPWR VGND sg13g2_decap_8
XFILLER_56_1000 VPWR VGND sg13g2_decap_8
X_14778_ _00579_ VGND VPWR _01302_ acc_sub.y\[7\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_90_196 VPWR VGND sg13g2_decap_8
XFILLER_90_185 VPWR VGND sg13g2_decap_8
XFILLER_17_794 VPWR VGND sg13g2_fill_2
XFILLER_32_720 VPWR VGND sg13g2_decap_8
X_13729_ VPWR _00280_ net67 VGND sg13g2_inv_1
X_07250_ _01583_ _01615_ _01614_ _01620_ VPWR VGND sg13g2_nand3_1
XFILLER_20_948 VPWR VGND sg13g2_decap_8
XFILLER_31_274 VPWR VGND sg13g2_fill_1
XFILLER_31_285 VPWR VGND sg13g2_decap_8
XFILLER_32_797 VPWR VGND sg13g2_decap_8
X_07181_ VGND VPWR _01547_ _01549_ _01553_ _01552_ sg13g2_a21oi_1
XFILLER_118_803 VPWR VGND sg13g2_decap_8
XFILLER_117_302 VPWR VGND sg13g2_fill_2
XFILLER_69_0 VPWR VGND sg13g2_decap_8
XFILLER_117_368 VPWR VGND sg13g2_fill_2
X_09822_ VPWR _03934_ acc_sum.y\[10\] VGND sg13g2_inv_1
XFILLER_87_937 VPWR VGND sg13g2_decap_8
X_09753_ net1664 _03868_ _03866_ _03869_ VPWR VGND sg13g2_nand3_1
XFILLER_100_235 VPWR VGND sg13g2_decap_4
X_08704_ net1817 acc_sum.add_renorm0.mantisa\[1\] _02917_ VPWR VGND sg13g2_nor2_1
XFILLER_58_149 VPWR VGND sg13g2_decap_8
XFILLER_39_341 VPWR VGND sg13g2_decap_8
XFILLER_95_981 VPWR VGND sg13g2_decap_8
X_09684_ VGND VPWR acc_sum.add_renorm0.exp\[1\] acc_sum.add_renorm0.exp\[0\] _03800_
+ acc_sum.add_renorm0.exp\[2\] sg13g2_a21oi_1
XFILLER_66_171 VPWR VGND sg13g2_fill_1
XFILLER_55_845 VPWR VGND sg13g2_fill_1
XFILLER_94_491 VPWR VGND sg13g2_fill_1
X_08635_ VPWR VGND _02856_ _02798_ _02855_ _02843_ _02857_ _02844_ sg13g2_a221oi_1
X_08566_ _02789_ _02733_ _02790_ VPWR VGND sg13g2_nor2_2
XFILLER_70_826 VPWR VGND sg13g2_fill_2
XFILLER_70_815 VPWR VGND sg13g2_decap_8
XFILLER_54_366 VPWR VGND sg13g2_decap_8
XFILLER_42_517 VPWR VGND sg13g2_decap_8
XFILLER_120_35 VPWR VGND sg13g2_decap_8
X_07517_ _01838_ VPWR _01839_ VGND acc_sub.exp_mant_logic0.b\[13\] _01837_ sg13g2_o21ai_1
Xfanout12 net13 net12 VPWR VGND sg13g2_buf_2
X_08497_ _02723_ net1708 fpdiv.divider0.remainder_reg\[4\] VPWR VGND sg13g2_nand2_1
Xfanout34 net39 net34 VPWR VGND sg13g2_buf_2
Xfanout23 net24 net23 VPWR VGND sg13g2_buf_2
Xfanout56 net71 net56 VPWR VGND sg13g2_buf_1
Xfanout45 net46 net45 VPWR VGND sg13g2_buf_1
X_07448_ _01775_ VPWR _01444_ VGND _01774_ net1748 sg13g2_o21ai_1
Xfanout89 net91 net89 VPWR VGND sg13g2_buf_2
Xfanout78 net80 net78 VPWR VGND sg13g2_buf_1
XFILLER_50_583 VPWR VGND sg13g2_fill_2
Xfanout67 net71 net67 VPWR VGND sg13g2_buf_1
XFILLER_11_959 VPWR VGND sg13g2_decap_8
XFILLER_22_274 VPWR VGND sg13g2_decap_8
XFILLER_109_814 VPWR VGND sg13g2_decap_8
X_07379_ _01728_ net1888 acc\[13\] VPWR VGND sg13g2_nand2_1
X_09118_ VGND VPWR _03203_ _03160_ _03299_ _03096_ sg13g2_a21oi_1
XFILLER_13_77 VPWR VGND sg13g2_decap_8
XFILLER_108_357 VPWR VGND sg13g2_fill_1
XFILLER_108_346 VPWR VGND sg13g2_fill_2
X_10390_ _04440_ _04438_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[5\] VPWR VGND sg13g2_nand2_1
X_09049_ _03235_ _03181_ net1791 VPWR VGND sg13g2_nand2_1
XFILLER_89_59 VPWR VGND sg13g2_decap_4
XFILLER_116_390 VPWR VGND sg13g2_fill_2
X_12060_ _05897_ _05889_ _05906_ VPWR VGND sg13g2_nor2_1
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_104_574 VPWR VGND sg13g2_fill_1
XFILLER_104_563 VPWR VGND sg13g2_decap_8
X_11011_ _04991_ VPWR _01104_ VGND net1813 _02802_ sg13g2_o21ai_1
XFILLER_77_414 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_89_285 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_46_801 VPWR VGND sg13g2_decap_8
XFILLER_38_63 VPWR VGND sg13g2_decap_8
X_12962_ _06733_ _06732_ net1961 VPWR VGND sg13g2_nand2_1
X_14701_ _00502_ VGND VPWR _01229_ acc_sum.y\[4\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_12893_ _06670_ net1717 _00012_ VPWR VGND sg13g2_nand2_1
XFILLER_73_653 VPWR VGND sg13g2_fill_2
XFILLER_73_642 VPWR VGND sg13g2_decap_8
XFILLER_61_804 VPWR VGND sg13g2_decap_8
X_11913_ net1881 fpmul.seg_reg0.q\[42\] _05786_ VPWR VGND sg13g2_nor2_1
XFILLER_45_344 VPWR VGND sg13g2_decap_8
XFILLER_72_152 VPWR VGND sg13g2_decap_8
XFILLER_45_388 VPWR VGND sg13g2_fill_1
X_14632_ _00433_ VGND VPWR _01164_ fp16_sum_pipe.add_renorm0.mantisa\[3\] clknet_leaf_108_clk
+ sg13g2_dfrbpq_2
X_11844_ VPWR _05742_ _05637_ VGND sg13g2_inv_1
XFILLER_127_1009 VPWR VGND sg13g2_decap_4
XFILLER_14_720 VPWR VGND sg13g2_fill_2
XFILLER_33_539 VPWR VGND sg13g2_fill_2
X_14563_ _00364_ VGND VPWR _01099_ acc_sum.seg_reg0.q\[26\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_11775_ _05672_ _05654_ _05678_ VPWR VGND sg13g2_and2_1
X_14494_ _00295_ VGND VPWR _01030_ fpdiv.divider0.divisor\[5\] clknet_leaf_85_clk
+ sg13g2_dfrbpq_1
X_13514_ VPWR _00065_ net37 VGND sg13g2_inv_1
XFILLER_14_786 VPWR VGND sg13g2_decap_8
X_10726_ VPWR _04739_ _04737_ VGND sg13g2_inv_1
X_13445_ _07101_ VPWR _00781_ VGND _06918_ net1751 sg13g2_o21ai_1
X_10657_ _04654_ _04658_ _04664_ _04670_ VPWR VGND sg13g2_nor3_2
XFILLER_127_611 VPWR VGND sg13g2_decap_8
Xclkload15 clknet_5_31__leaf_clk clkload15/X VPWR VGND sg13g2_buf_8
Xclkload26 VPWR clkload26/Y clknet_leaf_129_clk VGND sg13g2_inv_1
XFILLER_62_7 VPWR VGND sg13g2_decap_4
Xclkload59 clknet_leaf_126_clk clkload59/Y VPWR VGND sg13g2_inv_4
X_13376_ _07064_ VPWR _00813_ VGND _06339_ net1694 sg13g2_o21ai_1
Xclkload37 clkload37/Y clknet_leaf_13_clk VPWR VGND sg13g2_inv_2
Xclkload48 clknet_leaf_109_clk clkload48/Y VPWR VGND sg13g2_inv_4
XFILLER_6_941 VPWR VGND sg13g2_decap_8
X_10588_ _04607_ acc_sub.x2\[5\] net1934 VPWR VGND sg13g2_nand2_1
XFILLER_126_154 VPWR VGND sg13g2_decap_8
XFILLER_114_305 VPWR VGND sg13g2_decap_8
XFILLER_114_349 VPWR VGND sg13g2_fill_2
XFILLER_114_338 VPWR VGND sg13g2_fill_1
X_12258_ _06104_ _06103_ _06094_ VPWR VGND sg13g2_nand2b_1
XFILLER_123_883 VPWR VGND sg13g2_decap_8
X_11209_ _02951_ _05148_ _05175_ VPWR VGND sg13g2_nor2_1
X_12189_ _06035_ _06032_ _06034_ VPWR VGND sg13g2_nand2_1
XFILLER_68_469 VPWR VGND sg13g2_decap_4
XFILLER_56_609 VPWR VGND sg13g2_decap_4
XFILLER_23_1010 VPWR VGND sg13g2_decap_4
XFILLER_110_1013 VPWR VGND sg13g2_fill_1
XFILLER_110_588 VPWR VGND sg13g2_fill_1
XFILLER_95_277 VPWR VGND sg13g2_decap_4
XFILLER_95_91 VPWR VGND sg13g2_fill_1
XFILLER_76_480 VPWR VGND sg13g2_decap_8
XFILLER_64_642 VPWR VGND sg13g2_decap_4
XFILLER_48_193 VPWR VGND sg13g2_decap_8
X_08420_ _02654_ _02650_ VPWR VGND sg13g2_inv_2
XFILLER_92_995 VPWR VGND sg13g2_decap_8
XFILLER_64_664 VPWR VGND sg13g2_fill_1
XFILLER_37_889 VPWR VGND sg13g2_decap_8
XFILLER_24_506 VPWR VGND sg13g2_decap_8
XFILLER_63_196 VPWR VGND sg13g2_fill_2
XFILLER_17_591 VPWR VGND sg13g2_fill_2
XFILLER_24_539 VPWR VGND sg13g2_decap_8
X_08351_ VPWR _02594_ _02593_ VGND sg13g2_inv_1
X_07302_ _01668_ net1784 acc_sub.add_renorm0.mantisa\[6\] VPWR VGND sg13g2_nand2_1
X_08282_ _02529_ VPWR _02530_ VGND _02469_ _02322_ sg13g2_o21ai_1
XFILLER_20_734 VPWR VGND sg13g2_decap_8
X_07233_ _01604_ _01603_ _01542_ VPWR VGND sg13g2_nand2_1
Xclkload9 clknet_5_19__leaf_clk clkload9/X VPWR VGND sg13g2_buf_8
XFILLER_20_756 VPWR VGND sg13g2_decap_8
XFILLER_118_611 VPWR VGND sg13g2_fill_2
X_07164_ VPWR _01536_ _01535_ VGND sg13g2_inv_1
XFILLER_117_154 VPWR VGND sg13g2_decap_8
XFILLER_115_35 VPWR VGND sg13g2_decap_8
XFILLER_113_371 VPWR VGND sg13g2_decap_4
X_09805_ _03915_ _03918_ _03919_ VPWR VGND sg13g2_nor2b_1
X_07997_ _02264_ fp16_sum_pipe.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_inv_2
X_09736_ _03852_ _03851_ _03678_ VPWR VGND sg13g2_xnor2_1
XFILLER_101_588 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_27_311 VPWR VGND sg13g2_decap_8
XFILLER_55_653 VPWR VGND sg13g2_decap_8
X_08618_ VPWR _02840_ _02799_ VGND sg13g2_inv_1
XFILLER_83_995 VPWR VGND sg13g2_decap_8
XFILLER_28_889 VPWR VGND sg13g2_decap_8
X_09598_ _03711_ _03714_ _03715_ VPWR VGND sg13g2_nor2_1
XFILLER_42_325 VPWR VGND sg13g2_decap_8
X_08549_ VPWR _02773_ _02772_ VGND sg13g2_inv_1
XFILLER_24_21 VPWR VGND sg13g2_decap_8
XFILLER_11_712 VPWR VGND sg13g2_decap_8
X_11560_ _05442_ _05464_ _05465_ VPWR VGND sg13g2_nor2_2
X_10511_ VGND VPWR net1736 _04486_ _04554_ _04553_ sg13g2_a21oi_1
XFILLER_10_222 VPWR VGND sg13g2_decap_8
XFILLER_24_98 VPWR VGND sg13g2_decap_8
X_11491_ fpdiv.divider0.divisor\[5\] fp16_res_pipe.x2\[1\] net1944 _01030_ VPWR VGND
+ sg13g2_mux2_1
X_13230_ acc_sub.reg4en.q\[0\] _02576_ _06955_ VPWR VGND sg13g2_nor2_1
XFILLER_108_132 VPWR VGND sg13g2_fill_1
XFILLER_40_42 VPWR VGND sg13g2_decap_8
X_10442_ VGND VPWR _04488_ _04409_ _04491_ _04490_ sg13g2_a21oi_1
XFILLER_109_699 VPWR VGND sg13g2_fill_2
XFILLER_109_677 VPWR VGND sg13g2_fill_2
X_13161_ _06907_ _06901_ _06905_ VPWR VGND sg13g2_nand2_2
X_10373_ _04420_ _04422_ _04423_ VPWR VGND sg13g2_nor2_2
X_13092_ _06853_ VPWR _00886_ VGND fpmul.reg2en.q\[0\] _06655_ sg13g2_o21ai_1
X_12112_ VPWR _05958_ _05957_ VGND sg13g2_inv_1
XFILLER_123_168 VPWR VGND sg13g2_decap_8
X_12043_ _05889_ _05886_ _05888_ VPWR VGND sg13g2_nand2_1
XFILLER_3_966 VPWR VGND sg13g2_decap_8
XFILLER_2_465 VPWR VGND sg13g2_decap_8
XFILLER_120_820 VPWR VGND sg13g2_decap_8
XFILLER_104_382 VPWR VGND sg13g2_decap_8
XFILLER_78_756 VPWR VGND sg13g2_decap_8
XFILLER_66_918 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_120_897 VPWR VGND sg13g2_decap_8
XFILLER_59_970 VPWR VGND sg13g2_decap_4
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_46_653 VPWR VGND sg13g2_decap_4
X_13994_ VPWR _00545_ net9 VGND sg13g2_inv_1
XFILLER_18_344 VPWR VGND sg13g2_fill_2
XFILLER_80_409 VPWR VGND sg13g2_fill_1
X_12945_ acc\[2\] load_en _03983_ _06717_ VPWR VGND sg13g2_nand3_1
XFILLER_74_984 VPWR VGND sg13g2_fill_1
X_12876_ _06654_ _06650_ _06653_ _06499_ net1949 VPWR VGND sg13g2_a22oi_1
XFILLER_45_196 VPWR VGND sg13g2_decap_4
XFILLER_18_388 VPWR VGND sg13g2_fill_2
X_14615_ _00416_ VGND VPWR _01147_ fp16_sum_pipe.exp_mant_logic0.a\[10\] clknet_leaf_122_clk
+ sg13g2_dfrbpq_1
X_11827_ _05727_ _05496_ _05726_ _05724_ _05491_ VPWR VGND sg13g2_a22oi_1
XFILLER_33_347 VPWR VGND sg13g2_decap_4
X_14546_ _00347_ VGND VPWR _01082_ acc_sum.op_sign_logic0.mantisa_b\[9\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
XFILLER_14_561 VPWR VGND sg13g2_fill_2
X_11758_ VPWR _05662_ _05661_ VGND sg13g2_inv_1
X_10709_ _04647_ _04665_ _04722_ VPWR VGND sg13g2_nor2_1
Xclkload104 clkload104/Y clknet_leaf_61_clk VPWR VGND sg13g2_inv_2
X_14477_ _00278_ VGND VPWR _01015_ add_result\[2\] clknet_leaf_107_clk sg13g2_dfrbpq_1
X_11689_ VGND VPWR fp16_sum_pipe.add_renorm0.exp\[1\] fp16_sum_pipe.add_renorm0.exp\[0\]
+ _05593_ fp16_sum_pipe.add_renorm0.exp\[2\] sg13g2_a21oi_1
X_13428_ _07093_ net1720 instr\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_127_485 VPWR VGND sg13g2_decap_8
X_13359_ _07053_ VPWR _00819_ VGND _07018_ net1723 sg13g2_o21ai_1
Xplace1905 net1903 net1905 VPWR VGND sg13g2_buf_2
Xplace1916 net1913 net1916 VPWR VGND sg13g2_buf_1
Xplace1927 net1925 net1927 VPWR VGND sg13g2_buf_1
XFILLER_115_658 VPWR VGND sg13g2_decap_8
Xplace1938 fpdiv.reg1en.d\[0\] net1938 VPWR VGND sg13g2_buf_1
Xplace1949 net1948 net1949 VPWR VGND sg13g2_buf_2
XFILLER_5_270 VPWR VGND sg13g2_fill_2
XFILLER_114_168 VPWR VGND sg13g2_decap_8
X_07920_ fp16_sum_pipe.exp_mant_logic0.a\[11\] _02194_ _02195_ VPWR VGND sg13g2_nor2_1
XFILLER_111_831 VPWR VGND sg13g2_decap_8
XFILLER_69_745 VPWR VGND sg13g2_fill_2
XFILLER_110_330 VPWR VGND sg13g2_fill_1
X_07851_ _02146_ acc_sub.exp_mant_logic0.b\[0\] _01949_ acc_sub.exp_mant_logic0.b\[2\]
+ net1650 VPWR VGND sg13g2_a22oi_1
XFILLER_69_778 VPWR VGND sg13g2_decap_8
XFILLER_110_352 VPWR VGND sg13g2_fill_2
X_07782_ _02082_ net1649 net1794 VPWR VGND sg13g2_nand2_1
XFILLER_84_715 VPWR VGND sg13g2_decap_8
Xinput2 rst net2 VPWR VGND sg13g2_buf_1
XFILLER_56_428 VPWR VGND sg13g2_decap_8
XFILLER_56_406 VPWR VGND sg13g2_decap_8
XFILLER_110_396 VPWR VGND sg13g2_decap_8
X_09521_ VPWR _03638_ acc_sum.add_renorm0.mantisa\[8\] VGND sg13g2_inv_1
XFILLER_83_225 VPWR VGND sg13g2_decap_4
XFILLER_64_461 VPWR VGND sg13g2_decap_8
XFILLER_25_826 VPWR VGND sg13g2_fill_1
XFILLER_92_781 VPWR VGND sg13g2_decap_8
XFILLER_91_280 VPWR VGND sg13g2_fill_2
XFILLER_36_163 VPWR VGND sg13g2_decap_8
X_09452_ _03587_ net1832 fp16_res_pipe.seg_reg0.q\[23\] VPWR VGND sg13g2_nand2_1
X_08403_ VGND VPWR _02595_ _02638_ _02639_ _02603_ sg13g2_a21oi_1
XFILLER_52_678 VPWR VGND sg13g2_decap_8
X_09383_ _03530_ VPWR _03531_ VGND _03388_ _03529_ sg13g2_o21ai_1
XFILLER_24_369 VPWR VGND sg13g2_decap_4
X_08334_ _02574_ _02578_ _02579_ VPWR VGND sg13g2_nor2_1
XFILLER_20_542 VPWR VGND sg13g2_fill_1
X_08265_ _02515_ _02514_ _02475_ VPWR VGND sg13g2_nand2_1
XFILLER_20_564 VPWR VGND sg13g2_decap_4
X_07216_ _01582_ _01584_ _01587_ _01588_ VPWR VGND sg13g2_nor3_1
XFILLER_119_975 VPWR VGND sg13g2_decap_8
X_08196_ _02449_ _02451_ _02452_ _02453_ VPWR VGND sg13g2_nor3_1
XFILLER_118_485 VPWR VGND sg13g2_fill_1
XFILLER_118_463 VPWR VGND sg13g2_decap_4
X_07147_ VPWR _01519_ acc_sub.op_sign_logic0.mantisa_b\[7\] VGND sg13g2_inv_1
XFILLER_106_625 VPWR VGND sg13g2_decap_4
XFILLER_106_636 VPWR VGND sg13g2_fill_2
XFILLER_79_509 VPWR VGND sg13g2_fill_2
XFILLER_10_56 VPWR VGND sg13g2_decap_8
XFILLER_126_56 VPWR VGND sg13g2_decap_8
XFILLER_121_628 VPWR VGND sg13g2_fill_1
XFILLER_120_105 VPWR VGND sg13g2_decap_8
XFILLER_0_947 VPWR VGND sg13g2_decap_8
XFILLER_86_49 VPWR VGND sg13g2_fill_1
XFILLER_59_255 VPWR VGND sg13g2_fill_2
XFILLER_59_244 VPWR VGND sg13g2_fill_1
XFILLER_19_21 VPWR VGND sg13g2_decap_8
XFILLER_101_352 VPWR VGND sg13g2_decap_8
XFILLER_28_620 VPWR VGND sg13g2_fill_2
XFILLER_28_642 VPWR VGND sg13g2_decap_4
XFILLER_28_631 VPWR VGND sg13g2_fill_1
X_09719_ acc_sum.add_renorm0.exp\[4\] net1690 _03835_ VPWR VGND sg13g2_nor2_1
XFILLER_43_601 VPWR VGND sg13g2_decap_8
X_10991_ _04981_ VPWR _01114_ VGND net1933 _02210_ sg13g2_o21ai_1
X_12730_ _06534_ _06446_ _06529_ VPWR VGND sg13g2_xnor2_1
XFILLER_35_42 VPWR VGND sg13g2_decap_8
XFILLER_28_686 VPWR VGND sg13g2_fill_1
X_12661_ _06476_ _06468_ _06477_ VPWR VGND sg13g2_xor2_1
XFILLER_70_442 VPWR VGND sg13g2_fill_1
XFILLER_42_133 VPWR VGND sg13g2_decap_8
XFILLER_31_807 VPWR VGND sg13g2_fill_1
XFILLER_71_998 VPWR VGND sg13g2_fill_2
X_14400_ _00201_ VGND VPWR _00939_ div_result\[13\] clknet_leaf_89_clk sg13g2_dfrbpq_1
X_11612_ VPWR _05517_ _05415_ VGND sg13g2_inv_1
Xclkbuf_5_19__f_clk clknet_4_9_0_clk clknet_5_19__leaf_clk VPWR VGND sg13g2_buf_8
X_12592_ _06408_ _06395_ _06407_ VPWR VGND sg13g2_nand2_1
X_14331_ _00132_ VGND VPWR _00873_ piso.tx_bit_counter\[0\] clknet_leaf_56_clk sg13g2_dfrbpq_1
XFILLER_51_63 VPWR VGND sg13g2_decap_8
XFILLER_11_575 VPWR VGND sg13g2_fill_1
X_11543_ _05445_ _05447_ _05448_ VPWR VGND sg13g2_and2_1
X_11474_ _05388_ VPWR _01038_ VGND net1937 _05387_ sg13g2_o21ai_1
X_14262_ _00063_ VGND VPWR _00813_ acc_sub.x2\[11\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_51_74 VPWR VGND sg13g2_decap_8
X_14193_ VPWR _00744_ net91 VGND sg13g2_inv_1
X_13213_ VGND VPWR _06900_ sipo.receiving _06943_ net3 sg13g2_a21oi_1
X_10425_ _04474_ _04412_ _04416_ VPWR VGND sg13g2_nand2_2
XFILLER_125_956 VPWR VGND sg13g2_decap_8
X_13144_ _06887_ _06893_ _06886_ _00874_ VPWR VGND sg13g2_nor3_1
XFILLER_124_466 VPWR VGND sg13g2_fill_1
XFILLER_3_763 VPWR VGND sg13g2_decap_8
X_10356_ _04406_ _04404_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_112_639 VPWR VGND sg13g2_decap_4
XFILLER_97_328 VPWR VGND sg13g2_fill_1
X_13075_ _06817_ _06837_ _06842_ VPWR VGND _06841_ sg13g2_nand3b_1
X_10287_ _04352_ _04353_ _04355_ _04356_ VPWR VGND sg13g2_nor3_1
XFILLER_104_190 VPWR VGND sg13g2_decap_8
X_12026_ _05874_ _05842_ _05840_ VPWR VGND sg13g2_nand2_1
XFILLER_25_7 VPWR VGND sg13g2_decap_8
XFILLER_120_683 VPWR VGND sg13g2_decap_8
XFILLER_120_672 VPWR VGND sg13g2_fill_2
XFILLER_66_726 VPWR VGND sg13g2_decap_4
XFILLER_120_694 VPWR VGND sg13g2_fill_2
XFILLER_76_93 VPWR VGND sg13g2_decap_8
XFILLER_19_642 VPWR VGND sg13g2_fill_1
XFILLER_20_1013 VPWR VGND sg13g2_fill_1
XFILLER_62_910 VPWR VGND sg13g2_decap_8
X_13977_ VPWR _00528_ net16 VGND sg13g2_inv_1
XFILLER_19_664 VPWR VGND sg13g2_decap_8
X_12928_ _06702_ _06701_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_47_995 VPWR VGND sg13g2_decap_4
XFILLER_46_483 VPWR VGND sg13g2_fill_1
XFILLER_18_163 VPWR VGND sg13g2_decap_4
XFILLER_34_645 VPWR VGND sg13g2_decap_8
XFILLER_92_92 VPWR VGND sg13g2_decap_4
X_12859_ _00015_ net1730 net1701 _06638_ VPWR VGND sg13g2_nand3_1
XFILLER_14_380 VPWR VGND sg13g2_decap_8
X_14529_ _00330_ VGND VPWR _01065_ fpdiv.div_out\[4\] clknet_leaf_75_clk sg13g2_dfrbpq_2
XFILLER_30_862 VPWR VGND sg13g2_decap_4
XFILLER_119_238 VPWR VGND sg13g2_decap_8
X_08050_ _02316_ net1692 _02219_ VPWR VGND sg13g2_nand2b_1
XFILLER_116_912 VPWR VGND sg13g2_decap_8
Xplace1702 net1701 net1702 VPWR VGND sg13g2_buf_2
Xplace1735 net1734 net1735 VPWR VGND sg13g2_buf_2
Xplace1724 _07027_ net1724 VPWR VGND sg13g2_buf_2
Xplace1713 _06907_ net1713 VPWR VGND sg13g2_buf_2
XFILLER_51_0 VPWR VGND sg13g2_decap_8
XFILLER_116_989 VPWR VGND sg13g2_decap_8
XFILLER_115_455 VPWR VGND sg13g2_decap_8
Xplace1768 _03782_ net1768 VPWR VGND sg13g2_buf_2
XFILLER_89_829 VPWR VGND sg13g2_decap_8
Xplace1757 _05498_ net1757 VPWR VGND sg13g2_buf_1
Xplace1746 _04073_ net1746 VPWR VGND sg13g2_buf_2
X_08952_ VPWR _03138_ acc_sub.y\[14\] VGND sg13g2_inv_1
Xplace1779 _01779_ net1779 VPWR VGND sg13g2_buf_2
XFILLER_69_520 VPWR VGND sg13g2_decap_8
X_08883_ _03061_ _03062_ _03068_ _03070_ VPWR VGND sg13g2_nor3_2
X_07903_ _02178_ VPWR _01392_ VGND fp16_sum_pipe.reg1en.q\[0\] _02177_ sg13g2_o21ai_1
XFILLER_97_884 VPWR VGND sg13g2_fill_1
XFILLER_97_873 VPWR VGND sg13g2_decap_8
X_07834_ VPWR _02130_ acc_sub.exp_mant_logic0.b\[0\] VGND sg13g2_inv_1
XFILLER_38_951 VPWR VGND sg13g2_decap_4
XFILLER_112_14 VPWR VGND sg13g2_decap_8
X_07765_ _02067_ net1646 net1747 VPWR VGND sg13g2_nand2_1
XFILLER_65_770 VPWR VGND sg13g2_decap_8
XFILLER_38_973 VPWR VGND sg13g2_decap_8
XFILLER_37_461 VPWR VGND sg13g2_fill_1
X_07696_ _02002_ _02003_ _02004_ VPWR VGND sg13g2_nor2b_1
X_09504_ _03621_ acc_sum.add_renorm0.mantisa\[3\] acc_sum.add_renorm0.mantisa\[2\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_71_239 VPWR VGND sg13g2_fill_1
XFILLER_71_228 VPWR VGND sg13g2_decap_8
XFILLER_64_280 VPWR VGND sg13g2_decap_8
XFILLER_25_623 VPWR VGND sg13g2_decap_8
X_09435_ _03575_ VPWR _01264_ VGND net1834 _03574_ sg13g2_o21ai_1
XFILLER_24_177 VPWR VGND sg13g2_fill_2
XFILLER_52_497 VPWR VGND sg13g2_fill_1
X_09366_ _03437_ _03474_ _03516_ VPWR VGND sg13g2_nor2_1
XFILLER_12_328 VPWR VGND sg13g2_fill_1
XFILLER_12_339 VPWR VGND sg13g2_decap_8
X_08317_ VPWR _02562_ _02561_ VGND sg13g2_inv_1
X_09297_ _03443_ _03447_ _03450_ _03451_ VPWR VGND sg13g2_nor3_1
XFILLER_20_350 VPWR VGND sg13g2_decap_4
X_08248_ _02459_ _02340_ _02499_ VPWR VGND sg13g2_nor2_1
XFILLER_119_772 VPWR VGND sg13g2_decap_8
XFILLER_118_293 VPWR VGND sg13g2_decap_8
X_10210_ _04283_ _04284_ _04282_ _04285_ VPWR VGND sg13g2_nand3_1
X_08179_ _02434_ _02435_ _02436_ _02437_ VPWR VGND sg13g2_nor3_1
XFILLER_21_77 VPWR VGND sg13g2_fill_1
XFILLER_21_88 VPWR VGND sg13g2_decap_8
XFILLER_107_978 VPWR VGND sg13g2_decap_8
XFILLER_79_306 VPWR VGND sg13g2_decap_8
X_11190_ _05159_ net1809 net1680 acc_sum.op_sign_logic0.mantisa_a\[8\] net1759 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_122_959 VPWR VGND sg13g2_decap_8
XFILLER_106_488 VPWR VGND sg13g2_fill_1
X_10141_ _04128_ _04139_ net1662 _04222_ VPWR VGND sg13g2_nand3_1
XFILLER_88_862 VPWR VGND sg13g2_decap_8
XFILLER_43_1013 VPWR VGND sg13g2_fill_1
X_10072_ _04159_ net1643 net1746 VPWR VGND sg13g2_nand2_1
XFILLER_87_350 VPWR VGND sg13g2_decap_4
X_13900_ VPWR _00451_ net11 VGND sg13g2_inv_1
X_14880_ _00681_ VGND VPWR _01400_ acc_sub.exp_mant_logic0.b\[6\] clknet_leaf_58_clk
+ sg13g2_dfrbpq_2
XFILLER_90_515 VPWR VGND sg13g2_fill_1
XFILLER_63_707 VPWR VGND sg13g2_fill_2
X_13831_ VPWR _00382_ net51 VGND sg13g2_inv_1
XFILLER_29_962 VPWR VGND sg13g2_decap_8
X_13762_ VPWR _00313_ net129 VGND sg13g2_inv_1
XFILLER_56_770 VPWR VGND sg13g2_decap_8
X_10974_ net1835 fp16_res_pipe.y\[2\] _04974_ VPWR VGND sg13g2_nor2_1
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_44_921 VPWR VGND sg13g2_decap_4
XFILLER_15_100 VPWR VGND sg13g2_decap_8
XFILLER_16_612 VPWR VGND sg13g2_decap_8
X_12713_ _06519_ VPWR _00931_ VGND _06516_ net1741 sg13g2_o21ai_1
XFILLER_16_667 VPWR VGND sg13g2_fill_1
X_13693_ VPWR _00244_ net66 VGND sg13g2_inv_1
X_12644_ _06458_ _06459_ _06460_ VPWR VGND _06433_ sg13g2_nand3b_1
XFILLER_70_294 VPWR VGND sg13g2_fill_1
XFILLER_62_40 VPWR VGND sg13g2_decap_4
X_12575_ _06391_ fpdiv.reg_a_out\[11\] fpdiv.reg_b_out\[11\] VPWR VGND sg13g2_xnor2_1
XFILLER_12_862 VPWR VGND sg13g2_decap_8
XFILLER_30_158 VPWR VGND sg13g2_fill_2
X_14314_ _00115_ VGND VPWR _00857_ sipo.word\[2\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_11526_ fp16_sum_pipe.add_renorm0.mantisa\[2\] VPWR _05431_ VGND fp16_sum_pipe.add_renorm0.mantisa\[1\]
+ fp16_sum_pipe.add_renorm0.mantisa\[0\] sg13g2_o21ai_1
XFILLER_116_208 VPWR VGND sg13g2_decap_8
XFILLER_8_888 VPWR VGND sg13g2_decap_8
X_11457_ _05381_ acc_sub.x2\[2\] net1946 VPWR VGND sg13g2_nand2_1
X_14245_ _00046_ VGND VPWR _00796_ instr\[10\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_7_398 VPWR VGND sg13g2_decap_4
XFILLER_125_753 VPWR VGND sg13g2_decap_8
XFILLER_124_252 VPWR VGND sg13g2_decap_8
X_14176_ VPWR _00727_ net124 VGND sg13g2_inv_1
X_11388_ VPWR _05337_ fpdiv.div_out\[10\] VGND sg13g2_inv_1
X_10408_ VPWR _04458_ _04457_ VGND sg13g2_inv_1
XFILLER_97_125 VPWR VGND sg13g2_decap_4
X_13127_ net3 _06880_ VPWR VGND sg13g2_inv_4
X_10339_ VPWR _04389_ fp16_sum_pipe.seg_reg1.q\[20\] VGND sg13g2_inv_1
XFILLER_3_560 VPWR VGND sg13g2_decap_8
XFILLER_112_458 VPWR VGND sg13g2_decap_8
X_13058_ _05787_ _05789_ _06825_ _06826_ VPWR VGND _05791_ sg13g2_nand4_1
XFILLER_94_810 VPWR VGND sg13g2_fill_2
XFILLER_78_350 VPWR VGND sg13g2_fill_2
X_12009_ net1875 fpmul.seg_reg0.q\[22\] _05862_ VPWR VGND sg13g2_nor2_1
XFILLER_66_589 VPWR VGND sg13g2_decap_8
XFILLER_66_578 VPWR VGND sg13g2_fill_1
XFILLER_38_269 VPWR VGND sg13g2_fill_2
X_07550_ _01735_ _01737_ _01733_ _01865_ VPWR VGND _01739_ sg13g2_nand4_1
XFILLER_93_386 VPWR VGND sg13g2_decap_4
XFILLER_81_515 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_35_932 VPWR VGND sg13g2_decap_8
X_07481_ _01804_ acc_sub.exp_mant_logic0.b\[10\] VPWR VGND sg13g2_inv_2
X_09220_ VPWR _03374_ _03373_ VGND sg13g2_inv_1
XFILLER_99_0 VPWR VGND sg13g2_decap_8
XFILLER_50_957 VPWR VGND sg13g2_decap_4
X_09151_ VGND VPWR _03132_ net1800 _01297_ _03324_ sg13g2_a21oi_1
X_09082_ VGND VPWR _03248_ _03265_ _03266_ _03099_ sg13g2_a21oi_1
X_08102_ _02364_ _02365_ _02363_ _02366_ VPWR VGND sg13g2_nand3_1
X_08033_ _02298_ VPWR _02299_ VGND _02288_ net1692 sg13g2_o21ai_1
XFILLER_104_915 VPWR VGND sg13g2_decap_8
XFILLER_66_1013 VPWR VGND sg13g2_fill_1
XFILLER_116_786 VPWR VGND sg13g2_decap_8
XFILLER_115_252 VPWR VGND sg13g2_decap_8
XFILLER_107_69 VPWR VGND sg13g2_fill_1
XFILLER_103_436 VPWR VGND sg13g2_decap_8
XFILLER_88_147 VPWR VGND sg13g2_fill_1
X_09984_ _04070_ _04071_ _04069_ _04073_ VPWR VGND _04072_ sg13g2_nand4_1
X_08935_ _03121_ VPWR _03122_ VGND _02979_ _03092_ sg13g2_o21ai_1
XFILLER_69_372 VPWR VGND sg13g2_decap_8
XFILLER_123_35 VPWR VGND sg13g2_decap_8
X_08866_ VGND VPWR _03051_ _03052_ _03053_ net1785 sg13g2_a21oi_1
XFILLER_112_992 VPWR VGND sg13g2_decap_8
XFILLER_111_480 VPWR VGND sg13g2_decap_4
XFILLER_85_843 VPWR VGND sg13g2_fill_2
XFILLER_84_331 VPWR VGND sg13g2_fill_2
XFILLER_29_214 VPWR VGND sg13g2_decap_4
X_08797_ _01647_ _02982_ _02983_ _02984_ VPWR VGND sg13g2_nor3_1
X_07817_ _02112_ _02113_ _02111_ _02114_ VPWR VGND sg13g2_nand3_1
XFILLER_29_247 VPWR VGND sg13g2_decap_8
X_07748_ _02053_ _02052_ _01944_ VPWR VGND sg13g2_nand2_1
XFILLER_57_589 VPWR VGND sg13g2_fill_1
XFILLER_53_751 VPWR VGND sg13g2_fill_1
XFILLER_25_431 VPWR VGND sg13g2_decap_4
XFILLER_26_954 VPWR VGND sg13g2_decap_8
X_07679_ _01937_ _01933_ _01988_ VPWR VGND sg13g2_nor2_1
XFILLER_41_935 VPWR VGND sg13g2_decap_8
XFILLER_80_581 VPWR VGND sg13g2_decap_8
XFILLER_40_423 VPWR VGND sg13g2_decap_8
X_09418_ _03562_ _03407_ _03461_ VPWR VGND sg13g2_nand2b_1
X_10690_ _04703_ _04695_ _04679_ _04672_ net1710 VPWR VGND sg13g2_a22oi_1
XFILLER_25_497 VPWR VGND sg13g2_decap_8
X_09349_ _03361_ _03500_ _03501_ VPWR VGND sg13g2_nor2_2
XFILLER_32_21 VPWR VGND sg13g2_decap_8
X_12360_ VPWR _06206_ _06205_ VGND sg13g2_inv_1
X_11311_ _05268_ _05266_ _05267_ VPWR VGND sg13g2_nand2_1
XFILLER_5_803 VPWR VGND sg13g2_fill_2
XFILLER_107_731 VPWR VGND sg13g2_decap_8
X_12291_ _05939_ _05938_ _06136_ _06137_ VPWR VGND sg13g2_nand3_1
XFILLER_5_836 VPWR VGND sg13g2_decap_8
XFILLER_4_313 VPWR VGND sg13g2_decap_4
X_14030_ VPWR _00581_ net98 VGND sg13g2_inv_1
XFILLER_106_230 VPWR VGND sg13g2_fill_2
X_11242_ _05205_ VPWR _05206_ VGND _02957_ _05143_ sg13g2_o21ai_1
XFILLER_122_756 VPWR VGND sg13g2_decap_8
XFILLER_106_285 VPWR VGND sg13g2_fill_2
XFILLER_95_607 VPWR VGND sg13g2_decap_8
X_10124_ _04207_ fp16_res_pipe.exp_mant_logic0.a\[1\] net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[4\]
+ net1763 VPWR VGND sg13g2_a22oi_1
XFILLER_121_266 VPWR VGND sg13g2_decap_8
XFILLER_103_981 VPWR VGND sg13g2_decap_8
XFILLER_0_563 VPWR VGND sg13g2_fill_2
X_14932_ _00733_ VGND VPWR _01452_ acc_sub.exp_mant_logic0.a\[0\] clknet_leaf_56_clk
+ sg13g2_dfrbpq_2
XFILLER_48_523 VPWR VGND sg13g2_decap_8
XFILLER_48_512 VPWR VGND sg13g2_fill_2
X_10055_ VPWR _04143_ _04142_ VGND sg13g2_inv_1
XFILLER_63_504 VPWR VGND sg13g2_fill_1
XFILLER_48_578 VPWR VGND sg13g2_decap_8
X_14863_ _00664_ VGND VPWR _01387_ fp16_sum_pipe.seg_reg0.q\[25\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_1
XFILLER_91_846 VPWR VGND sg13g2_decap_8
X_13814_ VPWR _00365_ net75 VGND sg13g2_inv_1
XFILLER_36_729 VPWR VGND sg13g2_decap_8
XFILLER_90_345 VPWR VGND sg13g2_fill_1
X_14794_ _00595_ VGND VPWR _01318_ acc_sum.exp_mant_logic0.a\[7\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_44_751 VPWR VGND sg13g2_decap_8
XFILLER_17_954 VPWR VGND sg13g2_decap_8
XFILLER_28_280 VPWR VGND sg13g2_decap_8
X_13745_ VPWR _00296_ net118 VGND sg13g2_inv_1
X_10957_ _04962_ _04955_ _04865_ VPWR VGND sg13g2_nand2b_1
XFILLER_92_7 VPWR VGND sg13g2_decap_8
X_13676_ VPWR _00227_ net125 VGND sg13g2_inv_1
XFILLER_73_94 VPWR VGND sg13g2_decap_4
XFILLER_31_434 VPWR VGND sg13g2_fill_2
XFILLER_32_957 VPWR VGND sg13g2_decap_8
X_12627_ _06442_ _06423_ _06443_ VPWR VGND sg13g2_nor2_1
X_10888_ net1772 VPWR _04899_ VGND _04879_ _04898_ sg13g2_o21ai_1
XFILLER_117_517 VPWR VGND sg13g2_decap_8
X_12558_ _06374_ fpdiv.reg_a_out\[12\] fpdiv.reg_b_out\[12\] VPWR VGND sg13g2_xnor2_1
XFILLER_8_663 VPWR VGND sg13g2_decap_4
XFILLER_8_641 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_11_191 VPWR VGND sg13g2_decap_8
X_12489_ net1872 fpmul.seg_reg0.q\[6\] _06326_ VPWR VGND sg13g2_nor2_1
X_11509_ VPWR _05414_ _05413_ VGND sg13g2_inv_1
X_14228_ _00029_ VGND VPWR _00779_ sipo.shift_reg\[9\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_98_412 VPWR VGND sg13g2_decap_8
XFILLER_113_767 VPWR VGND sg13g2_decap_8
X_14159_ VPWR _00710_ net132 VGND sg13g2_inv_1
XFILLER_112_211 VPWR VGND sg13g2_fill_2
XFILLER_99_979 VPWR VGND sg13g2_decap_8
XFILLER_100_406 VPWR VGND sg13g2_decap_8
XFILLER_39_501 VPWR VGND sg13g2_decap_4
X_08720_ _02927_ net1819 acc_sum.seg_reg0.q\[25\] VPWR VGND sg13g2_nand2_1
XFILLER_79_692 VPWR VGND sg13g2_fill_1
XFILLER_94_651 VPWR VGND sg13g2_decap_8
X_08651_ VGND VPWR net1671 _02854_ _02871_ net1740 sg13g2_a21oi_1
XFILLER_78_191 VPWR VGND sg13g2_decap_8
XFILLER_67_887 VPWR VGND sg13g2_decap_8
XFILLER_66_342 VPWR VGND sg13g2_decap_4
XFILLER_39_556 VPWR VGND sg13g2_decap_8
XFILLER_14_0 VPWR VGND sg13g2_decap_8
X_07602_ _01829_ net1686 _01916_ VPWR VGND sg13g2_nor2_1
XFILLER_93_161 VPWR VGND sg13g2_decap_8
X_08582_ _02805_ VPWR _01347_ VGND net1814 _02729_ sg13g2_o21ai_1
XFILLER_82_879 VPWR VGND sg13g2_decap_8
XFILLER_81_334 VPWR VGND sg13g2_fill_2
XFILLER_54_559 VPWR VGND sg13g2_fill_2
XFILLER_54_548 VPWR VGND sg13g2_fill_2
XFILLER_26_239 VPWR VGND sg13g2_decap_8
X_07533_ _01853_ _01847_ acc_sub.exp_mant_logic0.a\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_81_378 VPWR VGND sg13g2_fill_2
X_07464_ VPWR _01787_ _01786_ VGND sg13g2_inv_1
XFILLER_50_743 VPWR VGND sg13g2_decap_4
XFILLER_50_721 VPWR VGND sg13g2_fill_2
XFILLER_34_294 VPWR VGND sg13g2_fill_1
X_09203_ _03358_ VPWR _01279_ VGND net1906 _03357_ sg13g2_o21ai_1
XFILLER_10_618 VPWR VGND sg13g2_fill_1
XFILLER_22_456 VPWR VGND sg13g2_fill_1
XFILLER_23_968 VPWR VGND sg13g2_decap_8
X_09134_ _03314_ _03135_ _03313_ VPWR VGND sg13g2_nand2_1
X_07395_ _01738_ VPWR _01460_ VGND net1895 _01737_ sg13g2_o21ai_1
X_09065_ VGND VPWR _03249_ _03199_ _03250_ _03099_ sg13g2_a21oi_1
XFILLER_118_35 VPWR VGND sg13g2_decap_8
X_08016_ _02280_ _02281_ _02282_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_828 VPWR VGND sg13g2_decap_8
XFILLER_89_467 VPWR VGND sg13g2_decap_8
XFILLER_77_607 VPWR VGND sg13g2_decap_4
XFILLER_58_810 VPWR VGND sg13g2_fill_2
X_09967_ _04060_ VPWR _01217_ VGND _04005_ _04054_ sg13g2_o21ai_1
X_08918_ _03105_ _02967_ _03007_ _02999_ _03004_ VPWR VGND sg13g2_a22oi_1
XFILLER_57_320 VPWR VGND sg13g2_decap_8
XFILLER_100_951 VPWR VGND sg13g2_decap_8
X_09898_ _03995_ fp16_res_pipe.exp_mant_logic0.b\[12\] VPWR VGND sg13g2_inv_2
XFILLER_18_707 VPWR VGND sg13g2_decap_8
X_08849_ VPWR _03036_ _03035_ VGND sg13g2_inv_1
XFILLER_57_375 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_73_868 VPWR VGND sg13g2_fill_2
X_11860_ VPWR _05757_ _05497_ VGND sg13g2_inv_1
X_11791_ _05608_ _05621_ _05642_ _05693_ VPWR VGND sg13g2_nand3_1
XFILLER_13_401 VPWR VGND sg13g2_decap_4
XFILLER_14_902 VPWR VGND sg13g2_decap_8
X_10811_ _04823_ _04775_ fp16_res_pipe.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_26_751 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_decap_8
X_13530_ VPWR _00081_ net34 VGND sg13g2_inv_1
X_10742_ _04753_ _04754_ _04755_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_272 VPWR VGND sg13g2_decap_4
XFILLER_43_42 VPWR VGND sg13g2_decap_8
XFILLER_13_445 VPWR VGND sg13g2_fill_2
XFILLER_14_979 VPWR VGND sg13g2_decap_8
X_13461_ _07110_ net1753 sipo.shift_reg\[3\] VPWR VGND sg13g2_nand2_1
X_10673_ _04685_ VPWR _04686_ VGND net1822 _04639_ sg13g2_o21ai_1
X_13392_ VGND VPWR _07010_ net1696 _00805_ _07072_ sg13g2_a21oi_1
X_12412_ _06257_ _06256_ _06258_ VPWR VGND sg13g2_xor2_1
XFILLER_127_848 VPWR VGND sg13g2_decap_8
XFILLER_126_336 VPWR VGND sg13g2_decap_8
X_12343_ _06189_ net1856 net1869 VPWR VGND sg13g2_nand2_1
XFILLER_5_600 VPWR VGND sg13g2_decap_8
X_12274_ _06120_ _06119_ _05965_ VPWR VGND sg13g2_nand2_1
X_14013_ VPWR _00564_ net75 VGND sg13g2_inv_1
X_11225_ _02957_ _05173_ _05190_ VPWR VGND sg13g2_nor2_1
XFILLER_4_154 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_122_564 VPWR VGND sg13g2_decap_8
X_11156_ _05126_ _05073_ _05124_ _05075_ net1808 VPWR VGND sg13g2_a22oi_1
XFILLER_1_850 VPWR VGND sg13g2_decap_8
XFILLER_110_759 VPWR VGND sg13g2_decap_8
X_11087_ _05062_ net1760 acc_sum.seg_reg0.q\[25\] VPWR VGND sg13g2_nand2_1
XFILLER_68_94 VPWR VGND sg13g2_fill_2
XFILLER_67_117 VPWR VGND sg13g2_decap_8
X_10107_ _04191_ net1642 net1746 VPWR VGND sg13g2_nand2_1
X_14915_ _00716_ VGND VPWR _01435_ acc_sub.seg_reg0.q\[25\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_76_662 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_decap_4
XFILLER_0_393 VPWR VGND sg13g2_decap_8
X_10038_ _04126_ _04124_ VPWR VGND sg13g2_inv_2
XFILLER_76_673 VPWR VGND sg13g2_fill_2
XFILLER_76_684 VPWR VGND sg13g2_fill_2
XFILLER_36_559 VPWR VGND sg13g2_decap_8
XFILLER_36_537 VPWR VGND sg13g2_decap_8
X_14846_ _00647_ VGND VPWR _01370_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[8\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
X_14777_ _00578_ VGND VPWR _01301_ acc_sub.y\[6\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_91_698 VPWR VGND sg13g2_decap_8
XFILLER_63_356 VPWR VGND sg13g2_decap_8
XFILLER_17_762 VPWR VGND sg13g2_fill_1
X_11989_ _05840_ _05842_ _05843_ VPWR VGND sg13g2_nor2_1
X_13728_ VPWR _00279_ net63 VGND sg13g2_inv_1
XFILLER_44_581 VPWR VGND sg13g2_fill_2
XFILLER_31_231 VPWR VGND sg13g2_fill_2
X_13659_ VPWR _00210_ net62 VGND sg13g2_inv_1
XFILLER_20_927 VPWR VGND sg13g2_decap_8
X_07180_ VPWR _01552_ _01551_ VGND sg13g2_inv_1
XFILLER_76_2 VPWR VGND sg13g2_fill_1
XFILLER_118_859 VPWR VGND sg13g2_decap_8
XFILLER_9_983 VPWR VGND sg13g2_decap_8
XFILLER_101_704 VPWR VGND sg13g2_decap_8
XFILLER_99_787 VPWR VGND sg13g2_fill_2
XFILLER_98_264 VPWR VGND sg13g2_fill_2
X_09821_ _01236_ _03932_ _03933_ VPWR VGND sg13g2_nand2_1
XFILLER_87_916 VPWR VGND sg13g2_decap_8
X_09752_ _03864_ _03867_ _03860_ _03868_ VPWR VGND sg13g2_nand3_1
XFILLER_98_286 VPWR VGND sg13g2_fill_1
XFILLER_58_128 VPWR VGND sg13g2_decap_8
XFILLER_100_258 VPWR VGND sg13g2_decap_8
XFILLER_95_960 VPWR VGND sg13g2_decap_8
X_08703_ _02916_ _02816_ _02915_ VPWR VGND sg13g2_xnor2_1
XFILLER_67_662 VPWR VGND sg13g2_fill_1
XFILLER_67_651 VPWR VGND sg13g2_decap_4
XFILLER_39_320 VPWR VGND sg13g2_decap_8
X_09683_ VPWR _03799_ _03798_ VGND sg13g2_inv_1
X_08634_ VGND VPWR _02732_ _02789_ _02856_ _02731_ sg13g2_a21oi_1
XFILLER_82_643 VPWR VGND sg13g2_decap_4
XFILLER_82_632 VPWR VGND sg13g2_decap_4
XFILLER_66_183 VPWR VGND sg13g2_fill_2
XFILLER_54_345 VPWR VGND sg13g2_decap_8
XFILLER_120_14 VPWR VGND sg13g2_decap_8
X_08565_ acc_sum.op_sign_logic0.mantisa_b\[8\] acc_sum.op_sign_logic0.mantisa_a\[8\]
+ _02789_ VPWR VGND sg13g2_nor2b_2
X_07516_ VGND VPWR _01837_ _01727_ _01838_ net1782 sg13g2_a21oi_1
XFILLER_81_186 VPWR VGND sg13g2_fill_1
XFILLER_23_732 VPWR VGND sg13g2_decap_8
Xfanout13 net14 net13 VPWR VGND sg13g2_buf_2
X_08496_ _02722_ fpdiv.divider0.dividend\[4\] VPWR VGND sg13g2_inv_2
Xfanout24 net39 net24 VPWR VGND sg13g2_buf_2
Xfanout35 net38 net35 VPWR VGND sg13g2_buf_2
XFILLER_22_231 VPWR VGND sg13g2_fill_2
XFILLER_23_776 VPWR VGND sg13g2_decap_8
Xfanout46 net47 net46 VPWR VGND sg13g2_buf_2
X_07447_ _01775_ net1750 fpdiv.divider0.divisor\[4\] VPWR VGND sg13g2_nand2_1
Xfanout79 net80 net79 VPWR VGND sg13g2_buf_2
Xfanout57 net60 net57 VPWR VGND sg13g2_buf_2
Xfanout68 net70 net68 VPWR VGND sg13g2_buf_2
XFILLER_50_562 VPWR VGND sg13g2_decap_8
XFILLER_11_938 VPWR VGND sg13g2_decap_8
XFILLER_22_253 VPWR VGND sg13g2_decap_8
X_07378_ _01727_ acc_sub.exp_mant_logic0.a\[13\] VPWR VGND sg13g2_inv_2
XFILLER_7_909 VPWR VGND sg13g2_decap_8
XFILLER_13_56 VPWR VGND sg13g2_decap_8
X_09117_ _03297_ VPWR _03298_ VGND _03173_ _02999_ sg13g2_o21ai_1
X_09048_ _03231_ _03233_ _03234_ VPWR VGND sg13g2_and2_1
XFILLER_89_38 VPWR VGND sg13g2_decap_8
XFILLER_123_339 VPWR VGND sg13g2_decap_8
X_11010_ _04991_ acc_sum.exp_mant_logic0.a\[15\] net1813 VPWR VGND sg13g2_nand2_1
XFILLER_78_916 VPWR VGND sg13g2_decap_8
XFILLER_89_275 VPWR VGND sg13g2_decap_4
XFILLER_78_949 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_93_919 VPWR VGND sg13g2_decap_8
XFILLER_38_42 VPWR VGND sg13g2_decap_8
XFILLER_79_1012 VPWR VGND sg13g2_fill_2
X_12961_ VPWR _06732_ fpmul.reg_p_out\[1\] VGND sg13g2_inv_1
XFILLER_45_301 VPWR VGND sg13g2_decap_8
X_14700_ _00501_ VGND VPWR _01228_ acc_sum.y\[3\] clknet_leaf_47_clk sg13g2_dfrbpq_1
X_12892_ _06669_ _06668_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_72_131 VPWR VGND sg13g2_decap_8
X_11912_ _05785_ fpmul.reg_a_out\[3\] VPWR VGND sg13g2_inv_2
XFILLER_46_868 VPWR VGND sg13g2_decap_4
XFILLER_45_323 VPWR VGND sg13g2_decap_4
XFILLER_18_537 VPWR VGND sg13g2_fill_2
XFILLER_18_548 VPWR VGND sg13g2_fill_2
X_11843_ _05741_ VPWR _01022_ VGND net1756 _05740_ sg13g2_o21ai_1
X_14631_ _00432_ VGND VPWR _01163_ fp16_sum_pipe.add_renorm0.mantisa\[2\] clknet_leaf_108_clk
+ sg13g2_dfrbpq_2
XFILLER_61_838 VPWR VGND sg13g2_decap_8
XFILLER_54_74 VPWR VGND sg13g2_decap_8
XFILLER_26_581 VPWR VGND sg13g2_decap_8
XFILLER_26_592 VPWR VGND sg13g2_fill_2
X_14562_ _00363_ VGND VPWR _01098_ acc_sum.seg_reg0.q\[25\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_54_96 VPWR VGND sg13g2_fill_2
X_11774_ _01027_ _05676_ _05677_ VPWR VGND sg13g2_nand2_1
XFILLER_41_551 VPWR VGND sg13g2_fill_1
XFILLER_41_540 VPWR VGND sg13g2_decap_8
X_14493_ _00294_ VGND VPWR _01029_ fpdiv.divider0.divisor\[4\] clknet_leaf_86_clk
+ sg13g2_dfrbpq_2
X_13513_ VPWR _00064_ net35 VGND sg13g2_inv_1
XFILLER_70_62 VPWR VGND sg13g2_fill_1
X_13444_ _07101_ net1751 sipo.shift_reg\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_6_920 VPWR VGND sg13g2_decap_8
XFILLER_10_982 VPWR VGND sg13g2_decap_8
Xclkload16 clknet_leaf_140_clk clkload16/Y VPWR VGND sg13g2_inv_4
XFILLER_126_133 VPWR VGND sg13g2_decap_8
Xclkload38 VPWR clkload38/Y clknet_leaf_16_clk VGND sg13g2_inv_1
X_13375_ _07064_ net1695 sipo.word\[11\] VPWR VGND sg13g2_nand2_1
Xclkload27 VPWR clkload27/Y clknet_leaf_131_clk VGND sg13g2_inv_1
Xclkload49 clknet_leaf_110_clk clkload49/Y VPWR VGND sg13g2_inv_4
X_10587_ _04606_ VPWR _01143_ VGND net1927 _02267_ sg13g2_o21ai_1
X_12326_ _06169_ _06171_ _06158_ _06172_ VPWR VGND sg13g2_nand3_1
XFILLER_55_7 VPWR VGND sg13g2_decap_8
XFILLER_6_997 VPWR VGND sg13g2_decap_8
X_12257_ _06103_ _06101_ _06102_ VPWR VGND sg13g2_nand2_1
XFILLER_5_485 VPWR VGND sg13g2_decap_8
XFILLER_123_862 VPWR VGND sg13g2_decap_8
XFILLER_96_702 VPWR VGND sg13g2_decap_8
X_11208_ _02955_ _05173_ _05174_ VPWR VGND sg13g2_nor2_1
X_12188_ _06034_ _06033_ net1855 VPWR VGND sg13g2_nand2_1
XFILLER_95_212 VPWR VGND sg13g2_decap_8
X_11139_ _05108_ VPWR _05109_ VGND _05021_ net1698 sg13g2_o21ai_1
XFILLER_37_868 VPWR VGND sg13g2_decap_8
XFILLER_36_323 VPWR VGND sg13g2_decap_8
X_14829_ _00630_ VGND VPWR _01353_ fpdiv.divider0.remainder_reg\[8\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_2
XFILLER_92_974 VPWR VGND sg13g2_decap_8
XFILLER_36_367 VPWR VGND sg13g2_decap_8
X_08350_ _02593_ instr\[1\] instr\[0\] VPWR VGND sg13g2_nand2_1
X_07301_ _01666_ VPWR _01667_ VGND _01527_ _01665_ sg13g2_o21ai_1
XFILLER_32_551 VPWR VGND sg13g2_fill_1
X_08281_ _02529_ _02338_ fp16_sum_pipe.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
X_07232_ _01602_ VPWR _01603_ VGND _01556_ _01554_ sg13g2_o21ai_1
X_07163_ _01532_ _01534_ _01535_ VPWR VGND sg13g2_nor2_2
XFILLER_118_634 VPWR VGND sg13g2_decap_4
XFILLER_30_1004 VPWR VGND sg13g2_decap_8
XFILLER_118_645 VPWR VGND sg13g2_decap_8
XFILLER_117_133 VPWR VGND sg13g2_decap_8
XFILLER_106_829 VPWR VGND sg13g2_fill_2
XFILLER_99_540 VPWR VGND sg13g2_fill_1
XFILLER_59_404 VPWR VGND sg13g2_decap_8
XFILLER_115_14 VPWR VGND sg13g2_decap_8
XFILLER_114_895 VPWR VGND sg13g2_decap_8
XFILLER_113_383 VPWR VGND sg13g2_decap_8
X_09804_ net1664 VPWR _03918_ VGND _03860_ _03917_ sg13g2_o21ai_1
XFILLER_86_223 VPWR VGND sg13g2_fill_1
XFILLER_113_394 VPWR VGND sg13g2_fill_2
XFILLER_86_256 VPWR VGND sg13g2_decap_4
X_07996_ _02261_ _02262_ _02260_ _02263_ VPWR VGND sg13g2_nand3_1
X_09735_ _03851_ _03849_ VPWR VGND sg13g2_inv_2
XFILLER_68_993 VPWR VGND sg13g2_decap_4
XFILLER_67_470 VPWR VGND sg13g2_fill_2
X_09666_ VGND VPWR _03782_ _03783_ _03781_ _03749_ sg13g2_a21oi_2
XFILLER_67_492 VPWR VGND sg13g2_fill_2
X_08617_ VGND VPWR _02803_ _02806_ _01346_ _02839_ sg13g2_a21oi_1
XFILLER_83_974 VPWR VGND sg13g2_decap_8
XFILLER_70_602 VPWR VGND sg13g2_decap_8
X_09597_ _03710_ _03713_ _03714_ VPWR VGND sg13g2_nor2_1
XFILLER_82_484 VPWR VGND sg13g2_decap_8
XFILLER_70_613 VPWR VGND sg13g2_fill_1
X_08548_ _02772_ _02770_ acc_sum.op_sign_logic0.mantisa_a\[4\] VPWR VGND sg13g2_nand2_1
X_08479_ _02709_ fpdiv.divider0.remainder_reg\[8\] net1708 net1748 fpdiv.divider0.dividend\[8\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_51_893 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_143_clk clknet_5_0__leaf_clk clknet_leaf_143_clk VPWR VGND sg13g2_buf_8
XFILLER_23_584 VPWR VGND sg13g2_fill_2
X_11490_ fpdiv.divider0.divisor\[6\] fp16_res_pipe.x2\[2\] net1945 _01031_ VPWR VGND
+ sg13g2_mux2_1
X_10510_ VGND VPWR _04550_ _04552_ _04553_ net1736 sg13g2_a21oi_1
XFILLER_24_77 VPWR VGND sg13g2_decap_8
XFILLER_109_623 VPWR VGND sg13g2_fill_1
XFILLER_7_739 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_10_267 VPWR VGND sg13g2_decap_8
X_10441_ VPWR _04490_ _04489_ VGND sg13g2_inv_1
XFILLER_109_634 VPWR VGND sg13g2_fill_1
XFILLER_40_21 VPWR VGND sg13g2_decap_8
XFILLER_10_278 VPWR VGND sg13g2_fill_1
XFILLER_124_615 VPWR VGND sg13g2_fill_1
XFILLER_108_166 VPWR VGND sg13g2_decap_8
X_13160_ _06906_ _06905_ net1 VPWR VGND sg13g2_nand2_1
X_10372_ VPWR _04422_ _04421_ VGND sg13g2_inv_1
X_13091_ _06807_ net1700 _06852_ _06853_ VPWR VGND sg13g2_nand3_1
X_12111_ _05957_ fpmul.reg_a_out\[6\] net1868 VPWR VGND sg13g2_nand2_1
XFILLER_40_98 VPWR VGND sg13g2_decap_8
XFILLER_3_945 VPWR VGND sg13g2_decap_8
XFILLER_123_147 VPWR VGND sg13g2_decap_8
XFILLER_111_309 VPWR VGND sg13g2_fill_1
XFILLER_105_851 VPWR VGND sg13g2_fill_1
X_12042_ _05883_ _05887_ _05882_ _05888_ VPWR VGND sg13g2_nand3_1
XFILLER_2_444 VPWR VGND sg13g2_decap_8
XFILLER_105_895 VPWR VGND sg13g2_decap_8
XFILLER_104_372 VPWR VGND sg13g2_decap_4
XFILLER_77_223 VPWR VGND sg13g2_fill_1
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_120_876 VPWR VGND sg13g2_decap_8
XFILLER_92_204 VPWR VGND sg13g2_decap_8
XFILLER_77_289 VPWR VGND sg13g2_decap_8
X_13993_ VPWR _00544_ net9 VGND sg13g2_inv_1
XFILLER_19_813 VPWR VGND sg13g2_fill_1
X_12944_ VGND VPWR net1936 add_result\[2\] _06716_ net1950 sg13g2_a21oi_1
XFILLER_46_632 VPWR VGND sg13g2_fill_1
XFILLER_19_846 VPWR VGND sg13g2_fill_2
XFILLER_74_974 VPWR VGND sg13g2_fill_2
XFILLER_65_84 VPWR VGND sg13g2_decap_4
XFILLER_61_602 VPWR VGND sg13g2_decap_4
X_12875_ _06652_ _06651_ net1922 _06653_ VPWR VGND sg13g2_a21o_2
XFILLER_61_646 VPWR VGND sg13g2_decap_8
XFILLER_45_175 VPWR VGND sg13g2_decap_8
XFILLER_27_890 VPWR VGND sg13g2_decap_8
X_14614_ _00415_ VGND VPWR _01146_ fp16_sum_pipe.exp_mant_logic0.a\[9\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_2
X_11826_ _05726_ _05725_ _05711_ VPWR VGND sg13g2_nand2_1
XFILLER_81_50 VPWR VGND sg13g2_decap_4
XFILLER_60_189 VPWR VGND sg13g2_decap_8
X_14545_ _00346_ VGND VPWR _01081_ acc_sum.op_sign_logic0.mantisa_b\[8\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
Xclkbuf_leaf_134_clk clknet_5_3__leaf_clk clknet_leaf_134_clk VPWR VGND sg13g2_buf_8
X_11757_ _05660_ VPWR _05661_ VGND net1838 _04591_ sg13g2_o21ai_1
XFILLER_119_409 VPWR VGND sg13g2_fill_1
X_10708_ _04721_ _04672_ _04720_ _04681_ _04694_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_595 VPWR VGND sg13g2_decap_4
X_14476_ _00277_ VGND VPWR _01014_ add_result\[1\] clknet_leaf_99_clk sg13g2_dfrbpq_1
X_11688_ _05592_ _05591_ VPWR VGND sg13g2_inv_2
Xclkload105 clknet_leaf_62_clk clkload105/X VPWR VGND sg13g2_buf_8
X_13427_ _07092_ VPWR _00790_ VGND _07006_ net1719 sg13g2_o21ai_1
X_10639_ _04652_ _04651_ fp16_res_pipe.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_2
X_13358_ _07053_ net1723 fp16_res_pipe.x2\[1\] VPWR VGND sg13g2_nand2_1
Xplace1906 net1902 net1906 VPWR VGND sg13g2_buf_2
XFILLER_6_750 VPWR VGND sg13g2_fill_1
Xplace1917 net1916 net1917 VPWR VGND sg13g2_buf_1
XFILLER_115_637 VPWR VGND sg13g2_decap_8
Xplace1939 net1938 net1939 VPWR VGND sg13g2_buf_1
X_12309_ _06155_ _06108_ _06084_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_260 VPWR VGND sg13g2_decap_4
Xplace1928 net1927 net1928 VPWR VGND sg13g2_buf_1
XFILLER_114_147 VPWR VGND sg13g2_decap_8
X_13289_ _07004_ acc_sub.y\[5\] net1711 acc_sum.y\[5\] net1728 VPWR VGND sg13g2_a22oi_1
XFILLER_111_810 VPWR VGND sg13g2_decap_8
XFILLER_96_521 VPWR VGND sg13g2_fill_1
XFILLER_96_510 VPWR VGND sg13g2_fill_2
X_07850_ _02141_ _02144_ _02145_ VPWR VGND sg13g2_nor2_1
XFILLER_96_554 VPWR VGND sg13g2_decap_4
XFILLER_69_768 VPWR VGND sg13g2_decap_4
XFILLER_111_887 VPWR VGND sg13g2_decap_8
X_07781_ _02081_ net1795 net1646 net1747 net1650 VPWR VGND sg13g2_a22oi_1
XFILLER_68_289 VPWR VGND sg13g2_decap_8
XFILLER_68_278 VPWR VGND sg13g2_decap_4
X_09520_ VPWR _03637_ _03624_ VGND sg13g2_inv_1
Xinput3 ss net3 VPWR VGND sg13g2_buf_2
XFILLER_92_760 VPWR VGND sg13g2_decap_8
XFILLER_65_974 VPWR VGND sg13g2_decap_8
XFILLER_64_495 VPWR VGND sg13g2_decap_8
XFILLER_52_635 VPWR VGND sg13g2_decap_8
X_09451_ _03586_ fp16_res_pipe.add_renorm0.exp\[1\] VPWR VGND sg13g2_inv_2
XFILLER_101_49 VPWR VGND sg13g2_decap_8
XFILLER_101_27 VPWR VGND sg13g2_fill_2
X_08402_ _02638_ _02563_ _02612_ VPWR VGND sg13g2_nand2_1
XFILLER_52_657 VPWR VGND sg13g2_decap_8
XFILLER_40_819 VPWR VGND sg13g2_fill_2
X_09382_ VGND VPWR _03529_ _03388_ _03530_ _03518_ sg13g2_a21oi_1
XFILLER_24_337 VPWR VGND sg13g2_fill_2
XFILLER_24_359 VPWR VGND sg13g2_fill_2
X_08333_ _02576_ _02578_ VPWR VGND sg13g2_inv_4
Xclkbuf_leaf_125_clk clknet_5_12__leaf_clk clknet_leaf_125_clk VPWR VGND sg13g2_buf_8
XFILLER_51_189 VPWR VGND sg13g2_decap_8
X_08264_ _02512_ _02513_ _02509_ _02514_ VPWR VGND sg13g2_nand3_1
XFILLER_32_381 VPWR VGND sg13g2_decap_8
XFILLER_20_576 VPWR VGND sg13g2_fill_2
X_07215_ _01587_ _01586_ _01547_ VPWR VGND sg13g2_nand2_1
XFILLER_119_954 VPWR VGND sg13g2_decap_8
XFILLER_118_431 VPWR VGND sg13g2_fill_1
XFILLER_69_1000 VPWR VGND sg13g2_fill_1
X_08195_ _02270_ net1648 _02452_ VPWR VGND sg13g2_nor2_1
X_07146_ acc_sub.op_sign_logic0.mantisa_b\[7\] _01517_ _01518_ VPWR VGND sg13g2_nor2_1
XFILLER_106_604 VPWR VGND sg13g2_fill_1
XFILLER_105_103 VPWR VGND sg13g2_decap_4
XFILLER_10_35 VPWR VGND sg13g2_decap_8
XFILLER_126_35 VPWR VGND sg13g2_decap_8
XFILLER_105_169 VPWR VGND sg13g2_decap_8
XFILLER_105_147 VPWR VGND sg13g2_fill_1
XFILLER_86_17 VPWR VGND sg13g2_decap_4
XFILLER_0_926 VPWR VGND sg13g2_decap_8
XFILLER_59_223 VPWR VGND sg13g2_decap_8
XFILLER_48_908 VPWR VGND sg13g2_fill_2
XFILLER_102_898 VPWR VGND sg13g2_decap_4
XFILLER_101_386 VPWR VGND sg13g2_decap_8
X_09718_ _03833_ VPWR _03834_ VGND _02924_ net1690 sg13g2_o21ai_1
XFILLER_74_248 VPWR VGND sg13g2_decap_4
X_10990_ _04981_ fp16_res_pipe.x2\[9\] net1932 VPWR VGND sg13g2_nand2_1
X_09649_ _03766_ _03655_ _03667_ _03684_ _03652_ VPWR VGND sg13g2_a22oi_1
XFILLER_70_421 VPWR VGND sg13g2_decap_8
XFILLER_43_613 VPWR VGND sg13g2_fill_1
XFILLER_42_112 VPWR VGND sg13g2_decap_8
XFILLER_35_21 VPWR VGND sg13g2_decap_8
XFILLER_15_315 VPWR VGND sg13g2_fill_1
XFILLER_16_827 VPWR VGND sg13g2_decap_8
XFILLER_28_698 VPWR VGND sg13g2_decap_8
X_12660_ _06476_ _06469_ _06475_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_668 VPWR VGND sg13g2_fill_1
XFILLER_70_487 VPWR VGND sg13g2_decap_8
XFILLER_35_98 VPWR VGND sg13g2_decap_8
X_11611_ _05481_ _05500_ _05515_ _05516_ VPWR VGND sg13g2_nor3_1
X_12591_ _06396_ _06406_ _06407_ VPWR VGND sg13g2_nor2b_1
X_14330_ _00131_ VGND VPWR _00872_ net4 clknet_leaf_81_clk sg13g2_dfrbpq_2
XFILLER_42_189 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_116_clk clknet_5_8__leaf_clk clknet_leaf_116_clk VPWR VGND sg13g2_buf_8
XFILLER_51_42 VPWR VGND sg13g2_decap_8
XFILLER_13_1010 VPWR VGND sg13g2_decap_4
X_11542_ _05447_ _05446_ _05436_ VPWR VGND sg13g2_nand2_1
X_11473_ _05388_ fp16_res_pipe.x2\[9\] net1940 VPWR VGND sg13g2_nand2_1
X_14261_ _00062_ VGND VPWR _00812_ acc_sub.x2\[10\] clknet_leaf_127_clk sg13g2_dfrbpq_2
X_14192_ VPWR _00743_ net90 VGND sg13g2_inv_1
X_13212_ VGND VPWR _06941_ net1714 _00855_ _06942_ sg13g2_a21oi_1
X_10424_ _04473_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[0\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[0\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_125_935 VPWR VGND sg13g2_decap_8
X_13143_ VGND VPWR _06882_ piso.tx_bit_counter\[0\] _06893_ piso.tx_bit_counter\[1\]
+ sg13g2_a21oi_1
XFILLER_97_307 VPWR VGND sg13g2_decap_8
XFILLER_3_742 VPWR VGND sg13g2_decap_8
X_10355_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[6\] _04404_ _04405_ VPWR VGND sg13g2_nor2_1
XFILLER_78_521 VPWR VGND sg13g2_decap_8
X_13074_ VGND VPWR _06819_ _06840_ _06841_ _06814_ sg13g2_a21oi_1
X_10286_ _04354_ _04233_ _04355_ VPWR VGND sg13g2_nor2_1
XFILLER_120_640 VPWR VGND sg13g2_fill_1
XFILLER_78_532 VPWR VGND sg13g2_fill_1
X_12025_ _05873_ fpmul.seg_reg0.q\[17\] VPWR VGND sg13g2_inv_2
XFILLER_120_651 VPWR VGND sg13g2_decap_8
XFILLER_93_502 VPWR VGND sg13g2_fill_2
XFILLER_66_738 VPWR VGND sg13g2_decap_8
XFILLER_65_204 VPWR VGND sg13g2_decap_8
XFILLER_18_7 VPWR VGND sg13g2_decap_8
XFILLER_19_632 VPWR VGND sg13g2_fill_1
XFILLER_47_963 VPWR VGND sg13g2_fill_1
X_13976_ VPWR _00527_ net17 VGND sg13g2_inv_1
XFILLER_18_142 VPWR VGND sg13g2_decap_8
X_12927_ _06700_ VPWR _06701_ VGND net1962 _06698_ sg13g2_o21ai_1
XFILLER_62_944 VPWR VGND sg13g2_decap_4
XFILLER_46_495 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
X_12858_ _06636_ _06637_ _06626_ _00904_ VPWR VGND sg13g2_nand3_1
XFILLER_62_988 VPWR VGND sg13g2_fill_1
X_11809_ _05710_ _05604_ _05599_ VPWR VGND sg13g2_xnor2_1
XFILLER_15_882 VPWR VGND sg13g2_decap_8
XFILLER_33_156 VPWR VGND sg13g2_fill_1
X_12789_ _06565_ _06559_ _06574_ VPWR VGND sg13g2_nor2_2
Xclkbuf_leaf_107_clk clknet_5_14__leaf_clk clknet_leaf_107_clk VPWR VGND sg13g2_buf_8
XFILLER_42_690 VPWR VGND sg13g2_decap_4
XFILLER_30_841 VPWR VGND sg13g2_decap_8
XFILLER_119_217 VPWR VGND sg13g2_decap_8
X_14528_ _00329_ VGND VPWR _01064_ fpdiv.div_out\[3\] clknet_leaf_72_clk sg13g2_dfrbpq_1
X_14459_ _00260_ VGND VPWR _00998_ fpmul.seg_reg0.q\[44\] clknet_leaf_99_clk sg13g2_dfrbpq_1
XFILLER_127_294 VPWR VGND sg13g2_decap_8
XFILLER_115_423 VPWR VGND sg13g2_fill_1
XFILLER_115_401 VPWR VGND sg13g2_decap_8
Xplace1714 net1713 net1714 VPWR VGND sg13g2_buf_2
Xplace1725 net1724 net1725 VPWR VGND sg13g2_buf_2
Xplace1703 _04029_ net1703 VPWR VGND sg13g2_buf_2
Xplace1736 _04386_ net1736 VPWR VGND sg13g2_buf_2
XFILLER_116_968 VPWR VGND sg13g2_decap_8
Xplace1747 _02058_ net1747 VPWR VGND sg13g2_buf_2
Xplace1769 _03740_ net1769 VPWR VGND sg13g2_buf_2
XFILLER_89_808 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_8
Xplace1758 net1757 net1758 VPWR VGND sg13g2_buf_2
X_08951_ _03137_ VPWR _01310_ VGND _01498_ _03136_ sg13g2_o21ai_1
XFILLER_102_128 VPWR VGND sg13g2_fill_1
XFILLER_97_852 VPWR VGND sg13g2_decap_8
XFILLER_69_543 VPWR VGND sg13g2_fill_1
X_07902_ _02178_ net1843 fp16_sum_pipe.exp_mant_logic0.b\[15\] VPWR VGND sg13g2_nand2_1
X_07833_ _02124_ _02125_ _02128_ _02129_ VPWR VGND sg13g2_nor3_1
XFILLER_96_340 VPWR VGND sg13g2_fill_2
XFILLER_69_565 VPWR VGND sg13g2_decap_4
XFILLER_111_695 VPWR VGND sg13g2_fill_2
XFILLER_111_684 VPWR VGND sg13g2_decap_8
Xclkbuf_5_25__f_clk clknet_4_12_0_clk clknet_5_25__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_29_429 VPWR VGND sg13g2_fill_1
X_07764_ _01419_ _02065_ _02066_ VPWR VGND sg13g2_nand2_1
XFILLER_84_557 VPWR VGND sg13g2_decap_8
XFILLER_72_708 VPWR VGND sg13g2_fill_1
XFILLER_56_259 VPWR VGND sg13g2_fill_2
XFILLER_2_91 VPWR VGND sg13g2_decap_8
X_09503_ VPWR _03620_ acc_sum.add_renorm0.mantisa\[6\] VGND sg13g2_inv_1
X_07695_ _02003_ net1793 _01975_ _01871_ acc_sub.exp_mant_logic0.a\[0\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_65_782 VPWR VGND sg13g2_decap_8
XFILLER_53_922 VPWR VGND sg13g2_fill_1
XFILLER_64_292 VPWR VGND sg13g2_decap_8
XFILLER_53_955 VPWR VGND sg13g2_fill_1
XFILLER_53_944 VPWR VGND sg13g2_decap_8
X_09434_ _03575_ net1833 fp16_res_pipe.seg_reg0.q\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_13_808 VPWR VGND sg13g2_decap_8
XFILLER_24_134 VPWR VGND sg13g2_decap_8
XFILLER_53_988 VPWR VGND sg13g2_decap_4
XFILLER_40_605 VPWR VGND sg13g2_fill_2
XFILLER_13_819 VPWR VGND sg13g2_fill_1
XFILLER_123_1002 VPWR VGND sg13g2_decap_8
X_09365_ _03515_ _03436_ _03514_ VPWR VGND sg13g2_xnor2_1
XFILLER_123_1013 VPWR VGND sg13g2_fill_1
X_08316_ state\[3\] state\[2\] _02561_ VPWR VGND sg13g2_nor2_1
X_09296_ _03450_ _03449_ _03411_ VPWR VGND sg13g2_nand2_1
XFILLER_21_874 VPWR VGND sg13g2_fill_1
XFILLER_122_7 VPWR VGND sg13g2_decap_8
X_08247_ _02466_ _02349_ _02498_ VPWR VGND sg13g2_nor2_1
XFILLER_20_384 VPWR VGND sg13g2_decap_4
XFILLER_21_896 VPWR VGND sg13g2_decap_8
XFILLER_119_751 VPWR VGND sg13g2_decap_8
XFILLER_107_957 VPWR VGND sg13g2_decap_8
XFILLER_106_401 VPWR VGND sg13g2_fill_2
XFILLER_4_539 VPWR VGND sg13g2_decap_4
X_08178_ _02262_ net1648 _02436_ VPWR VGND sg13g2_nor2_1
XFILLER_21_56 VPWR VGND sg13g2_decap_8
X_07129_ VPWR _01501_ acc_sub.op_sign_logic0.mantisa_b\[10\] VGND sg13g2_inv_1
XFILLER_106_456 VPWR VGND sg13g2_fill_2
XFILLER_122_938 VPWR VGND sg13g2_decap_8
XFILLER_0_712 VPWR VGND sg13g2_decap_4
X_10140_ _01205_ _04220_ _04221_ VPWR VGND sg13g2_nand2_1
XFILLER_121_459 VPWR VGND sg13g2_fill_2
X_10071_ VPWR _04158_ _04156_ VGND sg13g2_inv_1
XFILLER_88_896 VPWR VGND sg13g2_decap_4
XFILLER_87_373 VPWR VGND sg13g2_decap_8
XFILLER_75_513 VPWR VGND sg13g2_decap_8
XFILLER_0_778 VPWR VGND sg13g2_decap_4
XFILLER_101_183 VPWR VGND sg13g2_decap_8
XFILLER_87_395 VPWR VGND sg13g2_decap_8
XFILLER_87_384 VPWR VGND sg13g2_fill_1
XFILLER_75_535 VPWR VGND sg13g2_fill_1
XFILLER_75_524 VPWR VGND sg13g2_fill_1
XFILLER_47_237 VPWR VGND sg13g2_fill_1
XFILLER_29_941 VPWR VGND sg13g2_decap_8
XFILLER_75_568 VPWR VGND sg13g2_fill_1
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
X_13830_ VPWR _00381_ net51 VGND sg13g2_inv_1
X_13761_ VPWR _00312_ net129 VGND sg13g2_inv_1
XFILLER_90_527 VPWR VGND sg13g2_decap_8
XFILLER_16_624 VPWR VGND sg13g2_fill_1
X_10973_ VGND VPWR _04971_ net1821 _04973_ _04972_ sg13g2_a21oi_1
XFILLER_90_549 VPWR VGND sg13g2_fill_2
X_12712_ _06519_ _06513_ _06518_ VPWR VGND sg13g2_nand2b_1
XFILLER_55_292 VPWR VGND sg13g2_decap_8
XFILLER_15_112 VPWR VGND sg13g2_decap_8
X_13692_ VPWR _00243_ net66 VGND sg13g2_inv_1
XFILLER_43_476 VPWR VGND sg13g2_decap_8
X_12643_ _06459_ net1852 _06400_ VPWR VGND sg13g2_xnor2_1
XFILLER_62_52 VPWR VGND sg13g2_decap_8
XFILLER_30_126 VPWR VGND sg13g2_decap_4
XFILLER_31_649 VPWR VGND sg13g2_decap_4
X_12574_ fpdiv.reg_b_out\[10\] _05365_ _06390_ VPWR VGND sg13g2_nor2_1
XFILLER_12_841 VPWR VGND sg13g2_decap_8
X_14313_ _00114_ VGND VPWR _00856_ sipo.word\[1\] clknet_leaf_21_clk sg13g2_dfrbpq_2
XFILLER_7_14 VPWR VGND sg13g2_decap_8
X_11525_ VPWR _05430_ _05428_ VGND sg13g2_inv_1
X_14244_ _00045_ VGND VPWR _00795_ instr\[9\] clknet_leaf_16_clk sg13g2_dfrbpq_1
XFILLER_8_867 VPWR VGND sg13g2_decap_8
XFILLER_7_366 VPWR VGND sg13g2_decap_8
XFILLER_125_732 VPWR VGND sg13g2_decap_8
XFILLER_109_283 VPWR VGND sg13g2_fill_2
X_11456_ VPWR _05380_ fpdiv.divider0.dividend\[6\] VGND sg13g2_inv_1
XFILLER_124_231 VPWR VGND sg13g2_decap_8
X_14175_ VPWR _00726_ net124 VGND sg13g2_inv_1
X_11387_ _01073_ _05335_ _05336_ VPWR VGND sg13g2_nand2_1
X_10407_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[10\] _02457_ _04457_ VPWR VGND sg13g2_nor2_1
XFILLER_113_949 VPWR VGND sg13g2_decap_8
XFILLER_98_638 VPWR VGND sg13g2_decap_8
X_13126_ _06879_ VPWR _00878_ VGND net1862 _06743_ sg13g2_o21ai_1
X_10338_ VGND VPWR _04386_ net1844 _01174_ _04388_ sg13g2_a21oi_1
XFILLER_112_437 VPWR VGND sg13g2_fill_2
XFILLER_98_649 VPWR VGND sg13g2_decap_4
XFILLER_79_852 VPWR VGND sg13g2_decap_4
X_13057_ fpmul.seg_reg0.q\[45\] fpmul.seg_reg0.q\[44\] fpmul.seg_reg0.q\[43\] fpmul.seg_reg0.q\[42\]
+ _06825_ VPWR VGND sg13g2_nor4_1
XFILLER_3_594 VPWR VGND sg13g2_decap_8
X_12008_ _05861_ _05856_ _05853_ VPWR VGND sg13g2_xnor2_1
X_10269_ _04338_ VPWR _04339_ VGND _04288_ _04227_ sg13g2_o21ai_1
XFILLER_78_395 VPWR VGND sg13g2_fill_1
XFILLER_38_237 VPWR VGND sg13g2_decap_8
XFILLER_54_719 VPWR VGND sg13g2_decap_8
X_13959_ VPWR _00510_ net96 VGND sg13g2_inv_1
XFILLER_93_376 VPWR VGND sg13g2_decap_4
XFILLER_53_229 VPWR VGND sg13g2_fill_2
XFILLER_53_218 VPWR VGND sg13g2_decap_8
XFILLER_35_911 VPWR VGND sg13g2_decap_8
XFILLER_19_462 VPWR VGND sg13g2_fill_1
X_07480_ acc_sub.exp_mant_logic0.b\[10\] _01733_ _01803_ VPWR VGND sg13g2_nor2_1
XFILLER_19_495 VPWR VGND sg13g2_decap_4
XFILLER_35_988 VPWR VGND sg13g2_decap_8
XFILLER_50_936 VPWR VGND sg13g2_decap_8
XFILLER_34_498 VPWR VGND sg13g2_decap_4
XFILLER_21_126 VPWR VGND sg13g2_decap_8
X_09150_ net1800 acc_sub.y\[2\] _03324_ VPWR VGND sg13g2_nor2_1
X_09081_ _03265_ _03196_ _03183_ VPWR VGND sg13g2_nand2_1
X_08101_ _02365_ _02343_ _02273_ VPWR VGND sg13g2_nand2_1
X_08032_ _02298_ net1692 _02285_ VPWR VGND sg13g2_nand2_1
XFILLER_116_765 VPWR VGND sg13g2_decap_8
XFILLER_115_231 VPWR VGND sg13g2_decap_8
XFILLER_103_415 VPWR VGND sg13g2_decap_8
XFILLER_27_1009 VPWR VGND sg13g2_decap_4
X_09983_ fp16_res_pipe.exp_mant_logic0.a\[2\] fp16_res_pipe.exp_mant_logic0.a\[1\]
+ fp16_res_pipe.exp_mant_logic0.a\[0\] _04072_ VPWR VGND sg13g2_nor3_1
X_08934_ _03121_ _03010_ _03001_ VPWR VGND sg13g2_nand2_1
XFILLER_115_297 VPWR VGND sg13g2_fill_1
XFILLER_112_971 VPWR VGND sg13g2_decap_8
XFILLER_97_671 VPWR VGND sg13g2_fill_1
XFILLER_123_14 VPWR VGND sg13g2_decap_8
X_08865_ _03052_ _02999_ _03001_ VPWR VGND sg13g2_nand2_1
XFILLER_85_822 VPWR VGND sg13g2_fill_1
X_08796_ acc_sub.add_renorm0.mantisa\[5\] acc_sub.add_renorm0.mantisa\[4\] acc_sub.add_renorm0.mantisa\[6\]
+ _02983_ VPWR VGND acc_sub.add_renorm0.mantisa\[3\] sg13g2_nand4_1
X_07816_ _02113_ _01975_ net1795 VPWR VGND sg13g2_nand2_1
XFILLER_57_546 VPWR VGND sg13g2_decap_4
X_07747_ _02052_ _02046_ _02051_ VPWR VGND sg13g2_nand2_1
XFILLER_83_29 VPWR VGND sg13g2_fill_1
XFILLER_26_933 VPWR VGND sg13g2_decap_8
XFILLER_72_549 VPWR VGND sg13g2_decap_4
XFILLER_25_410 VPWR VGND sg13g2_decap_8
XFILLER_25_443 VPWR VGND sg13g2_decap_8
X_07678_ _01987_ _01949_ acc_sub.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_40_402 VPWR VGND sg13g2_decap_8
XFILLER_16_56 VPWR VGND sg13g2_decap_8
XFILLER_25_465 VPWR VGND sg13g2_fill_1
XFILLER_25_476 VPWR VGND sg13g2_decap_8
X_09417_ _03501_ VPWR _03561_ VGND _03407_ _03559_ sg13g2_o21ai_1
XFILLER_13_638 VPWR VGND sg13g2_decap_8
XFILLER_40_468 VPWR VGND sg13g2_decap_8
X_09348_ VPWR _03500_ _03364_ VGND sg13g2_inv_1
XFILLER_12_137 VPWR VGND sg13g2_fill_1
XFILLER_40_479 VPWR VGND sg13g2_fill_2
XFILLER_8_119 VPWR VGND sg13g2_decap_8
XFILLER_21_682 VPWR VGND sg13g2_fill_1
XFILLER_126_507 VPWR VGND sg13g2_decap_4
X_11310_ _05267_ net1811 net1656 net1697 acc_sum.exp_mant_logic0.b\[4\] VPWR VGND
+ sg13g2_a22oi_1
X_09279_ _03432_ VPWR _03433_ VGND _03391_ _03431_ sg13g2_o21ai_1
XFILLER_126_529 VPWR VGND sg13g2_fill_1
X_12290_ VPWR _06136_ _05973_ VGND sg13g2_inv_1
X_11241_ _05205_ net1655 acc_sum.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_4_358 VPWR VGND sg13g2_decap_8
XFILLER_122_702 VPWR VGND sg13g2_fill_2
XFILLER_79_104 VPWR VGND sg13g2_decap_8
X_11172_ net1663 _05140_ _05141_ VPWR VGND sg13g2_nor2b_2
XFILLER_122_735 VPWR VGND sg13g2_decap_8
X_10123_ _04206_ _04205_ _04150_ VPWR VGND sg13g2_nand2_1
XFILLER_121_245 VPWR VGND sg13g2_decap_8
XFILLER_103_960 VPWR VGND sg13g2_decap_8
XFILLER_88_671 VPWR VGND sg13g2_decap_4
X_14931_ _00732_ VGND VPWR _01451_ fpdiv.divider0.divisor_reg\[11\] clknet_leaf_70_clk
+ sg13g2_dfrbpq_1
XFILLER_102_481 VPWR VGND sg13g2_fill_1
XFILLER_94_129 VPWR VGND sg13g2_decap_8
XFILLER_87_181 VPWR VGND sg13g2_decap_8
X_10054_ _04011_ _04137_ _04142_ VPWR VGND sg13g2_nor2_1
XFILLER_76_866 VPWR VGND sg13g2_fill_1
XFILLER_57_96 VPWR VGND sg13g2_decap_8
XFILLER_36_708 VPWR VGND sg13g2_decap_8
X_14862_ _00663_ VGND VPWR _01386_ fp16_sum_pipe.seg_reg0.q\[24\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_1
XFILLER_91_825 VPWR VGND sg13g2_decap_8
X_13813_ VPWR _00364_ net75 VGND sg13g2_inv_1
XFILLER_63_527 VPWR VGND sg13g2_fill_2
XFILLER_35_229 VPWR VGND sg13g2_fill_2
XFILLER_29_771 VPWR VGND sg13g2_fill_2
XFILLER_113_91 VPWR VGND sg13g2_decap_8
XFILLER_91_869 VPWR VGND sg13g2_fill_2
X_14793_ _00594_ VGND VPWR _01317_ acc_sum.exp_mant_logic0.a\[6\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_17_933 VPWR VGND sg13g2_decap_8
X_13744_ VPWR _00295_ net117 VGND sg13g2_inv_1
X_10956_ _04961_ VPWR _01129_ VGND _04960_ _04771_ sg13g2_o21ai_1
XFILLER_16_465 VPWR VGND sg13g2_fill_1
X_13675_ VPWR _00226_ net125 VGND sg13g2_inv_1
X_10887_ _04878_ _04860_ _04898_ VPWR VGND sg13g2_and2_1
XFILLER_31_413 VPWR VGND sg13g2_decap_8
XFILLER_32_936 VPWR VGND sg13g2_decap_8
X_12626_ _06441_ VPWR _06442_ VGND net1852 fpdiv.div_out\[4\] sg13g2_o21ai_1
XFILLER_31_446 VPWR VGND sg13g2_fill_2
XFILLER_85_7 VPWR VGND sg13g2_decap_4
X_12557_ fpdiv.reg_b_out\[11\] _05363_ _06373_ VPWR VGND sg13g2_nor2_1
XFILLER_11_170 VPWR VGND sg13g2_decap_8
X_12488_ _06325_ _06242_ _06245_ VPWR VGND sg13g2_xnor2_1
X_11508_ _05413_ net1840 fp16_sum_pipe.add_renorm0.mantisa\[4\] VPWR VGND sg13g2_nand2_1
X_11439_ net1940 fpdiv.reg_a_out\[8\] _05369_ VPWR VGND sg13g2_nor2_1
X_14227_ _00028_ VGND VPWR _00778_ sipo.shift_reg\[8\] clknet_leaf_12_clk sg13g2_dfrbpq_1
XFILLER_125_584 VPWR VGND sg13g2_fill_2
X_14158_ VPWR _00709_ net134 VGND sg13g2_inv_1
XFILLER_99_958 VPWR VGND sg13g2_decap_8
XFILLER_98_92 VPWR VGND sg13g2_decap_8
X_13109_ _06802_ _06866_ _06864_ _06867_ VPWR VGND sg13g2_nand3_1
XFILLER_4_881 VPWR VGND sg13g2_decap_8
X_14089_ VPWR _00640_ net40 VGND sg13g2_inv_1
XFILLER_113_1012 VPWR VGND sg13g2_fill_2
XFILLER_66_321 VPWR VGND sg13g2_decap_8
XFILLER_39_524 VPWR VGND sg13g2_decap_8
X_08650_ VGND VPWR _02869_ net1816 _01344_ _02870_ sg13g2_a21oi_1
X_07601_ VGND VPWR _01883_ _01810_ _01915_ _01809_ sg13g2_a21oi_1
XFILLER_94_685 VPWR VGND sg13g2_decap_4
XFILLER_82_836 VPWR VGND sg13g2_fill_1
XFILLER_54_527 VPWR VGND sg13g2_decap_8
XFILLER_26_218 VPWR VGND sg13g2_decap_8
X_08581_ _02804_ VPWR _02805_ VGND acc_sum.op_sign_logic0.s_b _02800_ sg13g2_o21ai_1
XFILLER_82_858 VPWR VGND sg13g2_fill_1
XFILLER_81_346 VPWR VGND sg13g2_decap_4
X_07532_ _01852_ _01844_ acc_sub.exp_mant_logic0.b\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_81_357 VPWR VGND sg13g2_decap_8
X_07463_ _01783_ _01785_ _01786_ VPWR VGND sg13g2_nor2_1
XFILLER_23_947 VPWR VGND sg13g2_decap_8
X_09202_ _03358_ acc_sub.x2\[0\] net1906 VPWR VGND sg13g2_nand2_1
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
X_09133_ _03313_ _03310_ _03312_ _03307_ net1786 VPWR VGND sg13g2_a22oi_1
X_07394_ _01738_ net1893 acc\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_50_799 VPWR VGND sg13g2_decap_4
XFILLER_33_1013 VPWR VGND sg13g2_fill_1
XFILLER_31_991 VPWR VGND sg13g2_decap_8
XFILLER_118_14 VPWR VGND sg13g2_decap_8
X_09064_ _03249_ _03248_ _03153_ VPWR VGND sg13g2_nand2_1
XFILLER_108_529 VPWR VGND sg13g2_decap_8
X_08015_ VGND VPWR _02232_ _02211_ _02281_ _02206_ sg13g2_a21oi_1
XFILLER_2_807 VPWR VGND sg13g2_decap_8
XFILLER_104_768 VPWR VGND sg13g2_fill_1
XFILLER_103_245 VPWR VGND sg13g2_decap_8
XFILLER_77_619 VPWR VGND sg13g2_decap_8
XFILLER_76_107 VPWR VGND sg13g2_decap_8
X_09966_ _04060_ fp16_res_pipe.exp_mant_logic0.a\[11\] _04056_ net1765 fp16_res_pipe.seg_reg0.q\[26\]
+ VPWR VGND sg13g2_a22oi_1
X_08917_ _03054_ _03074_ _03046_ _03104_ VPWR VGND _03103_ sg13g2_nand4_1
XFILLER_100_930 VPWR VGND sg13g2_decap_8
XFILLER_58_833 VPWR VGND sg13g2_decap_8
X_09897_ fp16_res_pipe.exp_mant_logic0.b\[12\] _03593_ _03994_ VPWR VGND sg13g2_nor2_1
X_08848_ _03035_ _03032_ _03034_ VPWR VGND sg13g2_nand2_1
XFILLER_94_28 VPWR VGND sg13g2_decap_8
XFILLER_85_630 VPWR VGND sg13g2_fill_2
XFILLER_69_192 VPWR VGND sg13g2_decap_4
XFILLER_58_866 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_96_clk clknet_5_12__leaf_clk clknet_leaf_96_clk VPWR VGND sg13g2_buf_8
XFILLER_40_1006 VPWR VGND sg13g2_decap_8
X_08779_ _02966_ acc_sub.add_renorm0.mantisa\[3\] acc_sub.add_renorm0.mantisa\[2\]
+ VPWR VGND sg13g2_nand2_2
XFILLER_72_324 VPWR VGND sg13g2_decap_8
XFILLER_57_398 VPWR VGND sg13g2_fill_1
XFILLER_27_77 VPWR VGND sg13g2_decap_8
X_11790_ VGND VPWR _05642_ _05621_ _05692_ _05608_ sg13g2_a21oi_1
X_10810_ _04822_ _04809_ _04724_ VPWR VGND sg13g2_xnor2_1
XFILLER_53_582 VPWR VGND sg13g2_decap_4
XFILLER_43_21 VPWR VGND sg13g2_decap_8
XFILLER_14_958 VPWR VGND sg13g2_decap_8
X_10741_ net1822 VPWR _04754_ VGND _04642_ _04740_ sg13g2_o21ai_1
X_13460_ _07109_ VPWR _00774_ VGND _06933_ net1753 sg13g2_o21ai_1
X_12411_ _06257_ _06030_ _06032_ _06033_ net1855 VPWR VGND sg13g2_a22oi_1
XFILLER_43_98 VPWR VGND sg13g2_decap_8
XFILLER_41_788 VPWR VGND sg13g2_decap_8
XFILLER_40_287 VPWR VGND sg13g2_decap_8
XFILLER_40_254 VPWR VGND sg13g2_decap_4
X_10672_ net1822 VPWR _04685_ VGND _04668_ _04684_ sg13g2_o21ai_1
X_13391_ acc_sub.x2\[3\] net1696 _07072_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_20_clk clknet_5_18__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_127_827 VPWR VGND sg13g2_decap_8
XFILLER_126_315 VPWR VGND sg13g2_decap_8
X_12342_ _06179_ _06177_ _06174_ _06188_ VPWR VGND sg13g2_nand3_1
XFILLER_111_0 VPWR VGND sg13g2_decap_8
X_12273_ _05946_ _05945_ _06118_ _06119_ VPWR VGND sg13g2_nand3_1
XFILLER_5_634 VPWR VGND sg13g2_fill_2
XFILLER_4_133 VPWR VGND sg13g2_decap_8
XFILLER_107_551 VPWR VGND sg13g2_decap_8
X_11224_ _01089_ _05188_ _05189_ VPWR VGND sg13g2_nand2_1
X_14012_ VPWR _00563_ net75 VGND sg13g2_inv_1
XFILLER_122_521 VPWR VGND sg13g2_decap_8
XFILLER_96_906 VPWR VGND sg13g2_fill_1
XFILLER_95_427 VPWR VGND sg13g2_decap_8
X_11086_ _05061_ _05052_ acc_sum.exp_mant_logic0.a\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_49_833 VPWR VGND sg13g2_decap_8
XFILLER_0_372 VPWR VGND sg13g2_decap_8
X_10106_ _04190_ _04189_ VPWR VGND sg13g2_inv_2
X_14914_ _00715_ VGND VPWR _01434_ acc_sub.seg_reg0.q\[24\] clknet_leaf_45_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_87_clk clknet_5_24__leaf_clk clknet_leaf_87_clk VPWR VGND sg13g2_buf_8
XFILLER_91_600 VPWR VGND sg13g2_decap_8
XFILLER_75_151 VPWR VGND sg13g2_decap_8
X_14845_ _00646_ VGND VPWR _01369_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[7\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
XFILLER_1_1011 VPWR VGND sg13g2_fill_2
X_14776_ _00577_ VGND VPWR _01300_ acc_sub.y\[5\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_91_677 VPWR VGND sg13g2_decap_8
XFILLER_84_94 VPWR VGND sg13g2_decap_8
X_11988_ VPWR _05842_ _05841_ VGND sg13g2_inv_1
XFILLER_51_519 VPWR VGND sg13g2_decap_8
XFILLER_44_560 VPWR VGND sg13g2_decap_8
XFILLER_32_700 VPWR VGND sg13g2_fill_2
X_13727_ VPWR _00278_ net64 VGND sg13g2_inv_1
XFILLER_16_273 VPWR VGND sg13g2_decap_8
XFILLER_17_796 VPWR VGND sg13g2_fill_1
X_10939_ _04945_ VPWR _04946_ VGND _04824_ _04822_ sg13g2_o21ai_1
XFILLER_31_210 VPWR VGND sg13g2_decap_8
XFILLER_20_906 VPWR VGND sg13g2_decap_8
X_13658_ VPWR _00209_ net68 VGND sg13g2_inv_1
XFILLER_31_265 VPWR VGND sg13g2_decap_8
X_12609_ _06424_ VPWR _06425_ VGND fpdiv.div_out\[11\] _05350_ sg13g2_o21ai_1
X_13589_ VPWR _00140_ net121 VGND sg13g2_inv_1
Xclkbuf_leaf_11_clk clknet_5_1__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
XFILLER_9_962 VPWR VGND sg13g2_decap_8
XFILLER_118_838 VPWR VGND sg13g2_decap_8
XFILLER_117_337 VPWR VGND sg13g2_fill_1
XFILLER_8_483 VPWR VGND sg13g2_decap_8
XFILLER_99_722 VPWR VGND sg13g2_fill_1
XFILLER_98_232 VPWR VGND sg13g2_decap_8
X_09820_ _03933_ _03782_ acc_sum.y\[11\] VPWR VGND sg13g2_nand2_1
X_09751_ _03867_ _03832_ VPWR VGND sg13g2_inv_2
X_08702_ _02915_ _02913_ _02914_ _02817_ net1740 VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_78_clk clknet_5_26__leaf_clk clknet_leaf_78_clk VPWR VGND sg13g2_buf_8
XFILLER_104_38 VPWR VGND sg13g2_fill_2
X_09682_ _03797_ VPWR _03798_ VGND net1807 _02924_ sg13g2_o21ai_1
XFILLER_94_460 VPWR VGND sg13g2_decap_8
XFILLER_82_611 VPWR VGND sg13g2_decap_8
XFILLER_66_151 VPWR VGND sg13g2_fill_2
XFILLER_55_803 VPWR VGND sg13g2_decap_8
XFILLER_27_516 VPWR VGND sg13g2_fill_2
XFILLER_94_482 VPWR VGND sg13g2_decap_8
X_08633_ _02855_ _02854_ _02792_ VPWR VGND sg13g2_nand2_1
XFILLER_55_858 VPWR VGND sg13g2_fill_2
XFILLER_54_335 VPWR VGND sg13g2_decap_4
X_08564_ _02788_ _02732_ VPWR VGND sg13g2_inv_2
XFILLER_82_688 VPWR VGND sg13g2_decap_4
XFILLER_81_165 VPWR VGND sg13g2_decap_8
XFILLER_70_828 VPWR VGND sg13g2_fill_1
X_07515_ _01837_ _01833_ _01836_ VPWR VGND sg13g2_nand2_2
XFILLER_70_839 VPWR VGND sg13g2_decap_8
XFILLER_35_582 VPWR VGND sg13g2_fill_1
X_08495_ _02721_ VPWR _01350_ VGND net1705 _02720_ sg13g2_o21ai_1
Xfanout36 net38 net36 VPWR VGND sg13g2_buf_1
XFILLER_50_541 VPWR VGND sg13g2_decap_4
Xfanout25 net28 net25 VPWR VGND sg13g2_buf_2
XFILLER_23_744 VPWR VGND sg13g2_fill_2
Xfanout47 net72 net47 VPWR VGND sg13g2_buf_2
Xfanout14 net15 net14 VPWR VGND sg13g2_buf_2
X_07446_ VPWR _01774_ fpdiv.divider0.divisor_reg\[4\] VGND sg13g2_inv_1
Xfanout69 net70 net69 VPWR VGND sg13g2_buf_1
Xfanout58 net60 net58 VPWR VGND sg13g2_buf_1
XFILLER_11_917 VPWR VGND sg13g2_decap_8
X_07377_ _01726_ VPWR _01466_ VGND net1886 _01725_ sg13g2_o21ai_1
XFILLER_10_427 VPWR VGND sg13g2_decap_8
XFILLER_13_35 VPWR VGND sg13g2_decap_8
X_09116_ _03297_ _03173_ net1704 VPWR VGND sg13g2_nand2_1
XFILLER_109_849 VPWR VGND sg13g2_decap_8
XFILLER_108_315 VPWR VGND sg13g2_fill_2
X_09047_ net1791 _03184_ _03232_ _03233_ VPWR VGND sg13g2_a21o_1
XFILLER_108_348 VPWR VGND sg13g2_fill_1
XFILLER_2_615 VPWR VGND sg13g2_decap_8
XFILLER_117_893 VPWR VGND sg13g2_decap_8
XFILLER_2_626 VPWR VGND sg13g2_fill_2
XFILLER_104_543 VPWR VGND sg13g2_fill_1
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_104_598 VPWR VGND sg13g2_decap_8
X_09949_ fp16_res_pipe.exp_mant_logic0.b\[14\] _03589_ _04045_ VPWR VGND sg13g2_nor2_1
XFILLER_38_21 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_69_clk clknet_5_31__leaf_clk clknet_leaf_69_clk VPWR VGND sg13g2_buf_8
XFILLER_77_449 VPWR VGND sg13g2_fill_1
XFILLER_86_994 VPWR VGND sg13g2_decap_8
X_12960_ _06731_ _06727_ _06730_ _06536_ net1948 VPWR VGND sg13g2_a22oi_1
XFILLER_58_685 VPWR VGND sg13g2_decap_4
XFILLER_58_663 VPWR VGND sg13g2_decap_8
XFILLER_85_493 VPWR VGND sg13g2_decap_8
X_12891_ _06667_ VPWR _06668_ VGND net1962 _06665_ sg13g2_o21ai_1
X_11911_ VGND VPWR net1880 _05783_ _00997_ _05784_ sg13g2_a21oi_1
XFILLER_46_836 VPWR VGND sg13g2_decap_8
XFILLER_38_98 VPWR VGND sg13g2_decap_8
XFILLER_61_817 VPWR VGND sg13g2_decap_8
X_11842_ _05741_ net1756 add_result\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_45_379 VPWR VGND sg13g2_decap_8
X_14630_ _00431_ VGND VPWR _01162_ fp16_sum_pipe.add_renorm0.mantisa\[1\] clknet_leaf_109_clk
+ sg13g2_dfrbpq_1
X_14561_ _00362_ VGND VPWR _01097_ acc_sum.seg_reg0.q\[24\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_72_187 VPWR VGND sg13g2_fill_1
XFILLER_72_165 VPWR VGND sg13g2_fill_2
XFILLER_54_891 VPWR VGND sg13g2_fill_1
XFILLER_54_42 VPWR VGND sg13g2_decap_8
X_13512_ VPWR _00063_ net37 VGND sg13g2_inv_1
X_11773_ _05677_ _05573_ add_result\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_110_70 VPWR VGND sg13g2_decap_8
X_14492_ _00293_ VGND VPWR net1947 fpdiv.reg1en.q\[0\] clknet_leaf_73_clk sg13g2_dfrbpq_1
XFILLER_13_265 VPWR VGND sg13g2_fill_2
XFILLER_14_799 VPWR VGND sg13g2_fill_2
X_10724_ _04667_ _04736_ _04735_ _04737_ VPWR VGND sg13g2_nand3_1
X_13443_ _07100_ VPWR _00782_ VGND _06916_ net1751 sg13g2_o21ai_1
X_10655_ _04642_ _04667_ _04668_ VPWR VGND sg13g2_nor2_1
XFILLER_10_961 VPWR VGND sg13g2_decap_8
Xclkload17 clknet_leaf_143_clk clkload17/Y VPWR VGND sg13g2_inv_4
XFILLER_127_668 VPWR VGND sg13g2_fill_1
XFILLER_126_112 VPWR VGND sg13g2_decap_8
X_12325_ _06171_ _06170_ _06159_ VPWR VGND sg13g2_nand2_1
Xclkload39 VPWR clkload39/Y clknet_leaf_15_clk VGND sg13g2_inv_1
Xclkload28 clknet_leaf_134_clk clkload28/Y VPWR VGND sg13g2_inv_4
X_10586_ _04606_ acc_sub.x2\[6\] net1932 VPWR VGND sg13g2_nand2_1
XFILLER_127_679 VPWR VGND sg13g2_decap_8
XFILLER_6_976 VPWR VGND sg13g2_decap_8
XFILLER_5_464 VPWR VGND sg13g2_decap_8
XFILLER_126_189 VPWR VGND sg13g2_decap_8
XFILLER_123_841 VPWR VGND sg13g2_decap_8
X_12256_ _06097_ _06099_ _06096_ _06102_ VPWR VGND sg13g2_nand3_1
XFILLER_48_7 VPWR VGND sg13g2_decap_8
X_11207_ _05173_ net1655 VPWR VGND sg13g2_inv_2
XFILLER_68_405 VPWR VGND sg13g2_fill_2
X_12187_ VPWR _06033_ _05991_ VGND sg13g2_inv_1
XFILLER_122_373 VPWR VGND sg13g2_fill_1
XFILLER_122_362 VPWR VGND sg13g2_decap_8
XFILLER_110_524 VPWR VGND sg13g2_decap_8
X_11138_ _05108_ net1698 _05022_ VPWR VGND sg13g2_nand2b_1
XFILLER_68_438 VPWR VGND sg13g2_decap_8
XFILLER_122_395 VPWR VGND sg13g2_decap_8
Xclkbuf_5_6__f_clk clknet_4_3_0_clk clknet_5_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_49_652 VPWR VGND sg13g2_fill_1
XFILLER_49_641 VPWR VGND sg13g2_decap_8
XFILLER_110_1004 VPWR VGND sg13g2_decap_8
X_11069_ _05046_ _05042_ _05026_ VPWR VGND sg13g2_nand2_2
XFILLER_49_674 VPWR VGND sg13g2_fill_1
XFILLER_49_663 VPWR VGND sg13g2_decap_8
XFILLER_37_814 VPWR VGND sg13g2_fill_2
XFILLER_36_302 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_0_clk clknet_5_1__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
XFILLER_92_953 VPWR VGND sg13g2_decap_8
X_14828_ _00629_ VGND VPWR _01352_ fpdiv.divider0.remainder_reg\[7\] clknet_leaf_74_clk
+ sg13g2_dfrbpq_2
X_07300_ VGND VPWR _01665_ _01527_ _01666_ _01656_ sg13g2_a21oi_1
X_14759_ _00560_ VGND VPWR _01283_ acc_sum.exp_mant_logic0.b\[4\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_60_861 VPWR VGND sg13g2_decap_4
X_08280_ _01365_ _02527_ _02528_ VPWR VGND sg13g2_nand2_1
XFILLER_32_563 VPWR VGND sg13g2_decap_8
X_07231_ _01602_ _01601_ _01559_ VPWR VGND sg13g2_nand2_1
X_07162_ acc_sub.op_sign_logic0.mantisa_a\[5\] _01533_ _01534_ VPWR VGND sg13g2_nor2_1
XFILLER_118_613 VPWR VGND sg13g2_fill_1
XFILLER_74_0 VPWR VGND sg13g2_decap_8
XFILLER_117_112 VPWR VGND sg13g2_decap_8
XFILLER_105_318 VPWR VGND sg13g2_fill_2
XFILLER_117_189 VPWR VGND sg13g2_decap_8
XFILLER_114_874 VPWR VGND sg13g2_decap_8
XFILLER_5_91 VPWR VGND sg13g2_decap_8
X_09803_ _03906_ _03916_ _03917_ VPWR VGND sg13g2_nor2_1
XFILLER_101_535 VPWR VGND sg13g2_fill_1
XFILLER_87_758 VPWR VGND sg13g2_decap_8
XFILLER_75_909 VPWR VGND sg13g2_decap_8
XFILLER_68_950 VPWR VGND sg13g2_fill_1
XFILLER_59_449 VPWR VGND sg13g2_fill_2
X_07995_ _02262_ fp16_sum_pipe.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_inv_2
XFILLER_74_408 VPWR VGND sg13g2_decap_8
XFILLER_68_972 VPWR VGND sg13g2_decap_8
XFILLER_39_140 VPWR VGND sg13g2_decap_8
XFILLER_28_803 VPWR VGND sg13g2_fill_1
X_09665_ _03782_ acc_sum.reg3en.q\[0\] VPWR VGND sg13g2_inv_2
XFILLER_83_953 VPWR VGND sg13g2_decap_8
X_08616_ _02808_ _02838_ _02839_ VPWR VGND sg13g2_nor2_1
X_09596_ acc_sum.add_renorm0.mantisa\[1\] _03708_ _03712_ _03713_ VPWR VGND sg13g2_nor3_1
XFILLER_55_699 VPWR VGND sg13g2_fill_2
XFILLER_55_688 VPWR VGND sg13g2_decap_8
XFILLER_54_165 VPWR VGND sg13g2_decap_8
XFILLER_43_839 VPWR VGND sg13g2_decap_8
X_08547_ acc_sum.op_sign_logic0.mantisa_a\[4\] _02770_ _02771_ VPWR VGND sg13g2_nor2_2
XFILLER_35_390 VPWR VGND sg13g2_fill_2
X_08478_ _02707_ VPWR _02708_ VGND fpdiv.divider0.remainder_reg\[7\] net1647 sg13g2_o21ai_1
XFILLER_51_872 VPWR VGND sg13g2_fill_1
XFILLER_11_703 VPWR VGND sg13g2_fill_2
XFILLER_23_563 VPWR VGND sg13g2_fill_2
XFILLER_24_56 VPWR VGND sg13g2_decap_8
X_07429_ _01762_ VPWR _01450_ VGND _01760_ _01756_ sg13g2_o21ai_1
XFILLER_11_758 VPWR VGND sg13g2_decap_8
XFILLER_7_729 VPWR VGND sg13g2_decap_4
X_10440_ _04489_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[6\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[6\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_11_769 VPWR VGND sg13g2_fill_2
XFILLER_40_77 VPWR VGND sg13g2_decap_8
X_10371_ _04421_ _04419_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_123_126 VPWR VGND sg13g2_decap_8
X_13090_ _06805_ VPWR _06852_ VGND _06751_ _06851_ sg13g2_o21ai_1
X_12110_ _05956_ _05951_ _05955_ VPWR VGND sg13g2_nand2_1
XFILLER_3_924 VPWR VGND sg13g2_decap_8
XFILLER_2_423 VPWR VGND sg13g2_decap_8
XFILLER_78_703 VPWR VGND sg13g2_decap_4
X_12041_ VPWR _05887_ _05885_ VGND sg13g2_inv_1
XFILLER_46_1012 VPWR VGND sg13g2_fill_2
XFILLER_77_202 VPWR VGND sg13g2_fill_2
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_120_855 VPWR VGND sg13g2_decap_8
X_13992_ VPWR _00543_ net9 VGND sg13g2_inv_1
X_12943_ _00008_ net1731 net1702 _06715_ VPWR VGND sg13g2_nand3_1
XFILLER_74_953 VPWR VGND sg13g2_decap_8
XFILLER_74_931 VPWR VGND sg13g2_decap_8
XFILLER_46_622 VPWR VGND sg13g2_fill_2
XFILLER_46_611 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_18_302 VPWR VGND sg13g2_decap_8
XFILLER_65_52 VPWR VGND sg13g2_decap_4
XFILLER_45_154 VPWR VGND sg13g2_decap_8
XFILLER_18_357 VPWR VGND sg13g2_decap_8
X_12874_ _06652_ net1909 fp16_res_pipe.y\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_60_113 VPWR VGND sg13g2_decap_8
XFILLER_61_658 VPWR VGND sg13g2_decap_4
XFILLER_42_850 VPWR VGND sg13g2_decap_8
X_14613_ _00414_ VGND VPWR _01145_ fp16_sum_pipe.exp_mant_logic0.a\[8\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_2
X_11825_ _05725_ _05591_ _05620_ VPWR VGND sg13g2_nand2b_1
XFILLER_121_91 VPWR VGND sg13g2_decap_8
X_14544_ _00345_ VGND VPWR _01080_ acc_sum.op_sign_logic0.mantisa_b\[7\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
XFILLER_42_861 VPWR VGND sg13g2_fill_2
XFILLER_14_563 VPWR VGND sg13g2_fill_1
X_11756_ _05660_ _05594_ net1838 VPWR VGND sg13g2_nand2_1
X_14475_ _00276_ VGND VPWR _01013_ add_result\[0\] clknet_leaf_98_clk sg13g2_dfrbpq_1
XFILLER_41_371 VPWR VGND sg13g2_decap_4
X_10707_ _04647_ _04719_ _04665_ _04720_ VPWR VGND sg13g2_nor3_2
X_13426_ _07092_ net1719 instr\[4\] VPWR VGND sg13g2_nand2_1
X_11687_ VGND VPWR _05583_ _05589_ _05591_ _05590_ sg13g2_a21oi_1
Xclkload106 clknet_leaf_68_clk clkload106/Y VPWR VGND sg13g2_inv_4
X_10638_ VPWR _04651_ _04650_ VGND sg13g2_inv_1
XFILLER_127_465 VPWR VGND sg13g2_decap_4
Xplace1907 load_en net1907 VPWR VGND sg13g2_buf_2
X_13357_ _07052_ VPWR _00820_ VGND _07014_ net1724 sg13g2_o21ai_1
X_10569_ VGND VPWR _03327_ net1931 _01152_ _04597_ sg13g2_a21oi_1
Xplace1918 net1917 net1918 VPWR VGND sg13g2_buf_1
XFILLER_114_126 VPWR VGND sg13g2_decap_8
X_12308_ VPWR _06154_ _06077_ VGND sg13g2_inv_1
X_13288_ _07003_ sipo.word\[5\] VPWR VGND sg13g2_inv_2
XFILLER_5_272 VPWR VGND sg13g2_fill_1
Xplace1929 net1928 net1929 VPWR VGND sg13g2_buf_1
X_12239_ _06085_ _06078_ _06084_ VPWR VGND sg13g2_xnor2_1
XFILLER_5_283 VPWR VGND sg13g2_fill_2
XFILLER_123_693 VPWR VGND sg13g2_decap_8
XFILLER_111_866 VPWR VGND sg13g2_decap_8
XFILLER_68_235 VPWR VGND sg13g2_fill_1
XFILLER_68_224 VPWR VGND sg13g2_decap_8
XFILLER_60_1009 VPWR VGND sg13g2_decap_4
X_07780_ _01417_ _02079_ _02080_ VPWR VGND sg13g2_nand2_1
XFILLER_110_354 VPWR VGND sg13g2_fill_1
XFILLER_96_577 VPWR VGND sg13g2_decap_4
XFILLER_65_942 VPWR VGND sg13g2_fill_2
XFILLER_49_482 VPWR VGND sg13g2_decap_8
XFILLER_49_471 VPWR VGND sg13g2_fill_1
XFILLER_37_677 VPWR VGND sg13g2_fill_2
X_09450_ _03585_ VPWR _01259_ VGND net1832 _03584_ sg13g2_o21ai_1
XFILLER_91_271 VPWR VGND sg13g2_decap_4
XFILLER_80_923 VPWR VGND sg13g2_fill_1
X_08401_ _02637_ _02620_ _02624_ VPWR VGND sg13g2_nand2_1
XFILLER_51_102 VPWR VGND sg13g2_decap_4
XFILLER_36_198 VPWR VGND sg13g2_decap_4
X_09381_ _03528_ VPWR _03529_ VGND _03431_ net1674 sg13g2_o21ai_1
XFILLER_51_179 VPWR VGND sg13g2_fill_1
XFILLER_32_360 VPWR VGND sg13g2_decap_8
X_08263_ _02513_ fp16_sum_pipe.exp_mant_logic0.b\[3\] _02338_ _02275_ fp16_sum_pipe.exp_mant_logic0.b\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_07214_ VPWR _01586_ _01585_ VGND sg13g2_inv_1
XFILLER_119_933 VPWR VGND sg13g2_decap_8
X_08194_ _02261_ _02450_ _02451_ VPWR VGND sg13g2_nor2_1
XFILLER_118_454 VPWR VGND sg13g2_decap_4
X_07145_ VPWR _01517_ acc_sub.op_sign_logic0.mantisa_a\[7\] VGND sg13g2_inv_1
XFILLER_69_1012 VPWR VGND sg13g2_fill_2
XFILLER_106_638 VPWR VGND sg13g2_fill_1
XFILLER_10_14 VPWR VGND sg13g2_decap_8
XFILLER_126_14 VPWR VGND sg13g2_decap_8
XFILLER_0_905 VPWR VGND sg13g2_decap_8
XFILLER_99_360 VPWR VGND sg13g2_decap_8
XFILLER_87_555 VPWR VGND sg13g2_decap_8
XFILLER_87_533 VPWR VGND sg13g2_decap_4
XFILLER_75_717 VPWR VGND sg13g2_decap_8
XFILLER_59_257 VPWR VGND sg13g2_fill_1
XFILLER_19_56 VPWR VGND sg13g2_decap_8
X_09717_ _03833_ net1690 _03796_ VPWR VGND sg13g2_nand2_1
XFILLER_74_216 VPWR VGND sg13g2_decap_8
XFILLER_28_622 VPWR VGND sg13g2_fill_1
XFILLER_90_709 VPWR VGND sg13g2_decap_4
XFILLER_67_290 VPWR VGND sg13g2_decap_8
XFILLER_56_953 VPWR VGND sg13g2_fill_1
X_09648_ _03764_ VPWR _03765_ VGND net1802 _03759_ sg13g2_o21ai_1
XFILLER_83_772 VPWR VGND sg13g2_decap_8
XFILLER_76_1005 VPWR VGND sg13g2_decap_8
XFILLER_71_934 VPWR VGND sg13g2_fill_2
XFILLER_71_923 VPWR VGND sg13g2_decap_8
X_09579_ _03695_ VPWR _03696_ VGND net1806 _03634_ sg13g2_o21ai_1
X_12590_ _06404_ _06405_ _06406_ VPWR VGND sg13g2_nor2_1
XFILLER_35_77 VPWR VGND sg13g2_decap_8
X_11610_ _05514_ VPWR _05515_ VGND net1836 _05505_ sg13g2_o21ai_1
XFILLER_24_883 VPWR VGND sg13g2_decap_8
XFILLER_51_21 VPWR VGND sg13g2_decap_8
X_11541_ fp16_sum_pipe.add_renorm0.mantisa\[7\] fp16_sum_pipe.add_renorm0.mantisa\[6\]
+ _05427_ _05446_ VPWR VGND sg13g2_nand3_1
XFILLER_50_190 VPWR VGND sg13g2_decap_8
XFILLER_11_544 VPWR VGND sg13g2_decap_4
XFILLER_11_566 VPWR VGND sg13g2_decap_8
X_11472_ VPWR _05387_ fpdiv.reg_b_out\[9\] VGND sg13g2_inv_1
X_14260_ _00061_ VGND VPWR _00811_ acc_sub.x2\[9\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_7_537 VPWR VGND sg13g2_decap_4
XFILLER_125_914 VPWR VGND sg13g2_decap_8
X_14191_ VPWR _00742_ net102 VGND sg13g2_inv_1
X_13211_ sipo.shift_reg\[1\] net1714 _06942_ VPWR VGND sg13g2_nor2_1
X_10423_ VPWR _04472_ _04471_ VGND sg13g2_inv_1
X_13142_ _00875_ _06882_ _06892_ _06888_ _06568_ VPWR VGND sg13g2_a22oi_1
X_10354_ VPWR _04404_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[6\] VGND sg13g2_inv_1
XFILLER_124_435 VPWR VGND sg13g2_fill_2
XFILLER_83_1009 VPWR VGND sg13g2_decap_4
XFILLER_4_0 VPWR VGND sg13g2_decap_8
X_13073_ _06840_ _06748_ _06818_ VPWR VGND sg13g2_nand2b_1
X_10285_ VPWR _04354_ fp16_res_pipe.exp_mant_logic0.b\[1\] VGND sg13g2_inv_1
XFILLER_111_129 VPWR VGND sg13g2_fill_2
X_12024_ VGND VPWR _05871_ net1873 _00972_ _05872_ sg13g2_a21oi_1
XFILLER_2_286 VPWR VGND sg13g2_decap_8
XFILLER_2_297 VPWR VGND sg13g2_fill_1
XFILLER_76_51 VPWR VGND sg13g2_fill_1
XFILLER_38_419 VPWR VGND sg13g2_fill_1
XFILLER_78_599 VPWR VGND sg13g2_fill_2
XFILLER_76_84 VPWR VGND sg13g2_fill_2
XFILLER_59_791 VPWR VGND sg13g2_decap_8
XFILLER_47_931 VPWR VGND sg13g2_fill_1
XFILLER_19_611 VPWR VGND sg13g2_decap_4
XFILLER_20_1004 VPWR VGND sg13g2_decap_8
XFILLER_81_709 VPWR VGND sg13g2_decap_8
XFILLER_74_761 VPWR VGND sg13g2_decap_8
XFILLER_62_901 VPWR VGND sg13g2_fill_1
X_13975_ VPWR _00526_ net16 VGND sg13g2_inv_1
XFILLER_19_655 VPWR VGND sg13g2_decap_4
X_12926_ _06700_ _06699_ net1961 VPWR VGND sg13g2_nand2_1
XFILLER_34_614 VPWR VGND sg13g2_fill_1
XFILLER_18_176 VPWR VGND sg13g2_fill_1
XFILLER_92_50 VPWR VGND sg13g2_decap_8
X_12857_ _06637_ _06574_ _00015_ VPWR VGND sg13g2_nand2_1
XFILLER_33_113 VPWR VGND sg13g2_decap_8
XFILLER_61_488 VPWR VGND sg13g2_decap_8
X_11808_ _05708_ _05648_ _05707_ _05709_ VPWR VGND sg13g2_nand3_1
XFILLER_15_861 VPWR VGND sg13g2_decap_8
X_12788_ _06573_ _06567_ _06571_ VPWR VGND sg13g2_nand2_1
X_14527_ _00328_ VGND VPWR _01063_ fpdiv.div_out\[2\] clknet_leaf_72_clk sg13g2_dfrbpq_1
X_14458_ _00259_ VGND VPWR _00997_ fpmul.seg_reg0.q\[43\] clknet_leaf_99_clk sg13g2_dfrbpq_1
X_14389_ _00190_ VGND VPWR _00928_ div_result\[2\] clknet_leaf_83_clk sg13g2_dfrbpq_1
X_13409_ _07083_ net1721 instr\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_127_273 VPWR VGND sg13g2_decap_8
Xplace1704 _02979_ net1704 VPWR VGND sg13g2_buf_2
XFILLER_116_947 VPWR VGND sg13g2_decap_8
Xplace1726 net1725 net1726 VPWR VGND sg13g2_buf_2
Xplace1715 _06907_ net1715 VPWR VGND sg13g2_buf_1
Xplace1748 _01756_ net1748 VPWR VGND sg13g2_buf_2
Xplace1759 _04993_ net1759 VPWR VGND sg13g2_buf_2
Xplace1737 net1736 net1737 VPWR VGND sg13g2_buf_2
X_08950_ _03137_ net1773 acc_sub.y\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_124_991 VPWR VGND sg13g2_decap_8
X_08881_ _03067_ _03021_ _03065_ _03068_ VPWR VGND sg13g2_nand3_1
XFILLER_116_1010 VPWR VGND sg13g2_decap_4
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_07901_ VPWR _02177_ fp16_sum_pipe.op_sign_logic0.s_b VGND sg13g2_inv_1
XFILLER_111_663 VPWR VGND sg13g2_decap_8
X_07832_ _02128_ _02126_ _02127_ VPWR VGND sg13g2_nand2_1
XFILLER_97_897 VPWR VGND sg13g2_decap_4
XFILLER_69_588 VPWR VGND sg13g2_decap_8
XFILLER_57_717 VPWR VGND sg13g2_decap_8
XFILLER_84_514 VPWR VGND sg13g2_fill_1
XFILLER_2_70 VPWR VGND sg13g2_decap_8
X_07763_ _02066_ net1794 net1669 acc_sub.op_sign_logic0.mantisa_b\[9\] net1781 VPWR
+ VGND sg13g2_a22oi_1
X_09502_ VPWR _03619_ acc_sum.add_renorm0.mantisa\[9\] VGND sg13g2_inv_1
XFILLER_84_569 VPWR VGND sg13g2_decap_8
XFILLER_49_290 VPWR VGND sg13g2_fill_1
XFILLER_37_452 VPWR VGND sg13g2_fill_1
XFILLER_112_49 VPWR VGND sg13g2_decap_8
X_07694_ _02000_ _02001_ _01999_ _02002_ VPWR VGND sg13g2_nand3_1
XFILLER_25_603 VPWR VGND sg13g2_decap_8
XFILLER_53_967 VPWR VGND sg13g2_decap_8
XFILLER_52_422 VPWR VGND sg13g2_decap_8
X_09433_ VPWR _03574_ fp16_res_pipe.add_renorm0.exp\[7\] VGND sg13g2_inv_1
XFILLER_36_1011 VPWR VGND sg13g2_fill_2
X_09364_ _03513_ VPWR _03514_ VGND _03433_ net1674 sg13g2_o21ai_1
XFILLER_25_669 VPWR VGND sg13g2_decap_4
X_08315_ _02560_ state\[1\] state\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_21_820 VPWR VGND sg13g2_fill_1
XFILLER_24_179 VPWR VGND sg13g2_fill_1
X_09295_ VPWR _03449_ _03448_ VGND sg13g2_inv_1
XFILLER_21_853 VPWR VGND sg13g2_fill_2
XFILLER_119_730 VPWR VGND sg13g2_decap_8
X_08246_ _02468_ _02223_ _02497_ VPWR VGND sg13g2_nor2_1
X_08177_ _02269_ _02349_ _02435_ VPWR VGND sg13g2_nor2_1
XFILLER_21_35 VPWR VGND sg13g2_decap_8
XFILLER_118_273 VPWR VGND sg13g2_decap_4
X_07128_ acc_sub.op_sign_logic0.mantisa_b\[10\] _01499_ _01500_ VPWR VGND sg13g2_nor2_1
XFILLER_115_7 VPWR VGND sg13g2_decap_8
XFILLER_107_936 VPWR VGND sg13g2_decap_8
XFILLER_4_518 VPWR VGND sg13g2_decap_8
XFILLER_97_28 VPWR VGND sg13g2_decap_8
XFILLER_122_917 VPWR VGND sg13g2_decap_8
XFILLER_115_991 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_fill_2
XFILLER_48_717 VPWR VGND sg13g2_decap_4
XFILLER_0_757 VPWR VGND sg13g2_decap_8
XFILLER_101_162 VPWR VGND sg13g2_fill_1
XFILLER_101_151 VPWR VGND sg13g2_decap_8
XFILLER_29_920 VPWR VGND sg13g2_decap_8
XFILLER_90_506 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
X_13760_ VPWR _00311_ net117 VGND sg13g2_inv_1
X_10972_ net1821 _04756_ _04972_ VPWR VGND sg13g2_nor2_1
XFILLER_29_997 VPWR VGND sg13g2_decap_8
X_12711_ VGND VPWR _06517_ _06511_ _06518_ net1734 sg13g2_a21oi_1
XFILLER_46_98 VPWR VGND sg13g2_decap_8
X_13691_ VPWR _00242_ net65 VGND sg13g2_inv_1
XFILLER_16_647 VPWR VGND sg13g2_decap_8
XFILLER_16_658 VPWR VGND sg13g2_fill_2
X_12642_ VPWR _06458_ _06457_ VGND sg13g2_inv_1
XFILLER_71_764 VPWR VGND sg13g2_decap_8
XFILLER_70_241 VPWR VGND sg13g2_decap_4
XFILLER_62_20 VPWR VGND sg13g2_decap_8
XFILLER_15_168 VPWR VGND sg13g2_decap_8
X_12573_ _06389_ _06387_ _06388_ VPWR VGND sg13g2_nand2_1
X_14312_ _00113_ VGND VPWR _00855_ sipo.word\[0\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_8_846 VPWR VGND sg13g2_decap_8
XFILLER_11_363 VPWR VGND sg13g2_decap_4
XFILLER_11_374 VPWR VGND sg13g2_decap_4
XFILLER_12_897 VPWR VGND sg13g2_decap_8
X_11455_ _05379_ VPWR _01048_ VGND net1947 _05378_ sg13g2_o21ai_1
X_14243_ _00044_ VGND VPWR _00794_ instr\[8\] clknet_leaf_13_clk sg13g2_dfrbpq_1
Xclkbuf_5_31__f_clk clknet_4_15_0_clk clknet_5_31__leaf_clk VPWR VGND sg13g2_buf_8
X_10406_ VPWR VGND _04455_ _04396_ _04450_ _04392_ _04456_ _04397_ sg13g2_a221oi_1
XFILLER_124_210 VPWR VGND sg13g2_decap_8
X_14174_ VPWR _00725_ net137 VGND sg13g2_inv_1
X_11386_ _05336_ net1761 acc_sum.op_sign_logic0.mantisa_b\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_125_788 VPWR VGND sg13g2_decap_8
XFILLER_113_928 VPWR VGND sg13g2_decap_8
X_13125_ _06802_ net1700 _06877_ _06879_ VPWR VGND _06878_ sg13g2_nand4_1
X_10337_ fp16_sum_pipe.seg_reg1.q\[21\] net1844 _04388_ VPWR VGND sg13g2_nor2_1
XFILLER_124_287 VPWR VGND sg13g2_decap_8
X_13056_ _06824_ _06822_ _06823_ VPWR VGND sg13g2_nand2_1
X_10268_ _04338_ _04190_ fp16_res_pipe.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_30_7 VPWR VGND sg13g2_decap_8
XFILLER_94_812 VPWR VGND sg13g2_fill_1
XFILLER_78_352 VPWR VGND sg13g2_fill_1
X_12007_ VGND VPWR _05859_ net1875 _00977_ _05860_ sg13g2_a21oi_1
XFILLER_121_994 VPWR VGND sg13g2_decap_8
XFILLER_120_482 VPWR VGND sg13g2_decap_8
X_10199_ _01200_ _04274_ _04275_ VPWR VGND sg13g2_nand2_1
XFILLER_66_569 VPWR VGND sg13g2_decap_8
XFILLER_66_558 VPWR VGND sg13g2_decap_4
X_13958_ VPWR _00509_ net96 VGND sg13g2_inv_1
XFILLER_46_260 VPWR VGND sg13g2_decap_8
XFILLER_19_474 VPWR VGND sg13g2_decap_8
X_12909_ acc\[5\] net1908 net1767 _06684_ VPWR VGND sg13g2_nand3_1
XFILLER_35_967 VPWR VGND sg13g2_decap_8
XFILLER_62_786 VPWR VGND sg13g2_fill_2
XFILLER_61_252 VPWR VGND sg13g2_decap_8
XFILLER_50_915 VPWR VGND sg13g2_decap_8
XFILLER_34_466 VPWR VGND sg13g2_fill_2
X_13889_ VPWR _00440_ net49 VGND sg13g2_inv_1
XFILLER_22_606 VPWR VGND sg13g2_decap_8
XFILLER_62_797 VPWR VGND sg13g2_fill_1
XFILLER_21_105 VPWR VGND sg13g2_decap_4
XFILLER_22_628 VPWR VGND sg13g2_fill_1
XFILLER_14_190 VPWR VGND sg13g2_decap_8
X_09080_ _03089_ VPWR _03264_ VGND _03245_ _03263_ sg13g2_o21ai_1
X_08100_ _02364_ net1645 fp16_sum_pipe.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_30_661 VPWR VGND sg13g2_decap_8
XFILLER_30_672 VPWR VGND sg13g2_fill_1
X_08031_ _02296_ _02196_ _02297_ VPWR VGND sg13g2_xor2_1
XFILLER_116_700 VPWR VGND sg13g2_fill_2
XFILLER_116_744 VPWR VGND sg13g2_decap_8
XFILLER_115_210 VPWR VGND sg13g2_decap_8
XFILLER_89_617 VPWR VGND sg13g2_fill_1
XFILLER_89_606 VPWR VGND sg13g2_decap_8
XFILLER_88_105 VPWR VGND sg13g2_decap_8
X_09982_ fp16_res_pipe.exp_mant_logic0.a\[6\] fp16_res_pipe.exp_mant_logic0.a\[5\]
+ fp16_res_pipe.exp_mant_logic0.a\[4\] fp16_res_pipe.exp_mant_logic0.a\[3\] _04071_
+ VPWR VGND sg13g2_nor4_1
X_08933_ _03120_ _03119_ VPWR VGND sg13g2_inv_2
XFILLER_88_116 VPWR VGND sg13g2_fill_2
XFILLER_112_950 VPWR VGND sg13g2_decap_8
XFILLER_97_661 VPWR VGND sg13g2_decap_4
XFILLER_97_650 VPWR VGND sg13g2_fill_2
X_08864_ VPWR VGND _02967_ _03050_ _03017_ _03014_ _03051_ _03004_ sg13g2_a221oi_1
XFILLER_85_845 VPWR VGND sg13g2_fill_1
X_08795_ _02982_ acc_sub.add_renorm0.mantisa\[7\] VPWR VGND sg13g2_inv_2
X_07815_ _02112_ _01989_ net1794 VPWR VGND sg13g2_nand2_1
XFILLER_84_333 VPWR VGND sg13g2_fill_1
X_07746_ _02047_ _02049_ _02050_ _02051_ VPWR VGND sg13g2_nor3_1
XFILLER_84_366 VPWR VGND sg13g2_decap_8
XFILLER_44_208 VPWR VGND sg13g2_fill_2
XFILLER_26_912 VPWR VGND sg13g2_decap_8
XFILLER_72_539 VPWR VGND sg13g2_fill_2
XFILLER_16_35 VPWR VGND sg13g2_decap_8
X_07677_ _01426_ _01985_ _01986_ VPWR VGND sg13g2_nand2_1
X_09416_ _03559_ _03407_ _03560_ VPWR VGND sg13g2_and2_1
XFILLER_26_989 VPWR VGND sg13g2_decap_8
XFILLER_52_285 VPWR VGND sg13g2_decap_8
XFILLER_52_274 VPWR VGND sg13g2_decap_8
XFILLER_12_105 VPWR VGND sg13g2_decap_8
XFILLER_12_127 VPWR VGND sg13g2_decap_4
XFILLER_13_628 VPWR VGND sg13g2_decap_4
XFILLER_16_79 VPWR VGND sg13g2_decap_4
XFILLER_52_296 VPWR VGND sg13g2_fill_1
X_09347_ _03498_ VPWR _03499_ VGND _03445_ _03497_ sg13g2_o21ai_1
X_09278_ VGND VPWR _03382_ _03385_ _03432_ _03379_ sg13g2_a21oi_1
XFILLER_32_56 VPWR VGND sg13g2_decap_8
X_08229_ _02483_ net1638 _02482_ VPWR VGND sg13g2_nand2_1
XFILLER_10_1003 VPWR VGND sg13g2_decap_8
XFILLER_106_232 VPWR VGND sg13g2_fill_1
XFILLER_106_210 VPWR VGND sg13g2_fill_1
X_11240_ _05203_ VPWR _05204_ VGND _02963_ _05026_ sg13g2_o21ai_1
XFILLER_4_337 VPWR VGND sg13g2_decap_8
XFILLER_122_714 VPWR VGND sg13g2_decap_8
XFILLER_106_254 VPWR VGND sg13g2_decap_8
X_11171_ _05139_ _05122_ _05140_ VPWR VGND sg13g2_nor2_1
XFILLER_121_224 VPWR VGND sg13g2_decap_8
X_10122_ _04205_ _04200_ _04204_ VPWR VGND sg13g2_nand2_1
XFILLER_88_650 VPWR VGND sg13g2_decap_8
XFILLER_79_149 VPWR VGND sg13g2_fill_2
XFILLER_0_565 VPWR VGND sg13g2_fill_1
X_14930_ _00731_ VGND VPWR _01450_ fpdiv.divider0.divisor_reg\[10\] clknet_leaf_70_clk
+ sg13g2_dfrbpq_1
XFILLER_88_694 VPWR VGND sg13g2_decap_8
XFILLER_87_160 VPWR VGND sg13g2_decap_8
XFILLER_48_503 VPWR VGND sg13g2_fill_1
XFILLER_0_598 VPWR VGND sg13g2_decap_4
XFILLER_87_193 VPWR VGND sg13g2_decap_4
XFILLER_75_322 VPWR VGND sg13g2_decap_8
XFILLER_48_558 VPWR VGND sg13g2_decap_4
X_14861_ _00662_ VGND VPWR _01385_ fp16_sum_pipe.seg_reg0.q\[23\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_1
X_13812_ VPWR _00363_ net78 VGND sg13g2_inv_1
XFILLER_35_219 VPWR VGND sg13g2_fill_2
XFILLER_17_912 VPWR VGND sg13g2_decap_8
XFILLER_113_70 VPWR VGND sg13g2_decap_8
X_14792_ _00593_ VGND VPWR _01316_ acc_sum.exp_mant_logic0.a\[5\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_13743_ VPWR _00294_ net118 VGND sg13g2_inv_1
XFILLER_44_775 VPWR VGND sg13g2_decap_8
X_10955_ _04961_ _04772_ fp16_res_pipe.y\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_17_989 VPWR VGND sg13g2_decap_8
XFILLER_32_915 VPWR VGND sg13g2_decap_8
X_13674_ VPWR _00225_ net125 VGND sg13g2_inv_1
XFILLER_44_786 VPWR VGND sg13g2_fill_1
X_10886_ _04897_ _04771_ VPWR VGND sg13g2_inv_2
XFILLER_31_403 VPWR VGND sg13g2_fill_1
X_12625_ _06441_ _05345_ net1852 VPWR VGND sg13g2_nand2_1
XFILLER_43_296 VPWR VGND sg13g2_decap_4
XFILLER_31_436 VPWR VGND sg13g2_fill_1
XFILLER_8_621 VPWR VGND sg13g2_decap_8
XFILLER_78_7 VPWR VGND sg13g2_decap_4
XFILLER_40_992 VPWR VGND sg13g2_decap_8
X_11507_ _05412_ _05411_ VPWR VGND sg13g2_inv_2
X_12487_ VGND VPWR _06323_ net1872 _00961_ _06324_ sg13g2_a21oi_1
XFILLER_8_698 VPWR VGND sg13g2_decap_8
X_11438_ VGND VPWR _05367_ net1937 _01054_ _05368_ sg13g2_a21oi_1
X_14226_ _00027_ VGND VPWR _00777_ sipo.shift_reg\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_1
X_14157_ VPWR _00708_ net130 VGND sg13g2_inv_1
XFILLER_99_937 VPWR VGND sg13g2_decap_8
X_11369_ _05319_ VPWR _05320_ VGND _03351_ _05183_ sg13g2_o21ai_1
XFILLER_4_860 VPWR VGND sg13g2_decap_8
X_13108_ _06866_ _06801_ _06865_ VPWR VGND sg13g2_nand2b_1
XFILLER_86_609 VPWR VGND sg13g2_decap_4
XFILLER_3_392 VPWR VGND sg13g2_decap_8
X_14088_ VPWR _00639_ net40 VGND sg13g2_inv_1
XFILLER_26_1010 VPWR VGND sg13g2_decap_4
XFILLER_79_683 VPWR VGND sg13g2_decap_8
X_13039_ VPWR _06807_ _06806_ VGND sg13g2_inv_1
XFILLER_121_791 VPWR VGND sg13g2_decap_8
XFILLER_94_642 VPWR VGND sg13g2_decap_4
XFILLER_39_536 VPWR VGND sg13g2_fill_2
X_07600_ VPWR _01914_ _01913_ VGND sg13g2_inv_1
X_08580_ VGND VPWR _02800_ _02802_ _02804_ _02803_ sg13g2_a21oi_1
XFILLER_66_388 VPWR VGND sg13g2_decap_8
X_07531_ _01850_ _01851_ _01846_ _01437_ VPWR VGND sg13g2_nand3_1
XFILLER_35_742 VPWR VGND sg13g2_decap_8
XFILLER_62_550 VPWR VGND sg13g2_decap_8
XFILLER_35_775 VPWR VGND sg13g2_decap_8
XFILLER_35_764 VPWR VGND sg13g2_fill_2
X_07462_ acc_sub.exp_mant_logic0.a\[13\] _01784_ _01785_ VPWR VGND sg13g2_nor2_1
XFILLER_50_723 VPWR VGND sg13g2_fill_1
XFILLER_23_926 VPWR VGND sg13g2_decap_8
X_07393_ VPWR _01737_ acc_sub.exp_mant_logic0.a\[8\] VGND sg13g2_inv_1
X_09201_ _03357_ acc_sum.exp_mant_logic0.b\[0\] VPWR VGND sg13g2_inv_2
X_09132_ _03089_ _03311_ _03166_ _03312_ VPWR VGND sg13g2_nand3_1
XFILLER_50_778 VPWR VGND sg13g2_decap_8
XFILLER_31_970 VPWR VGND sg13g2_decap_8
XFILLER_30_480 VPWR VGND sg13g2_decap_4
X_09063_ VPWR _03248_ _03197_ VGND sg13g2_inv_1
XFILLER_8_91 VPWR VGND sg13g2_decap_8
X_08014_ _02213_ _02279_ _02280_ VPWR VGND sg13g2_nor2_1
XFILLER_116_563 VPWR VGND sg13g2_fill_2
XFILLER_104_736 VPWR VGND sg13g2_decap_8
XFILLER_89_425 VPWR VGND sg13g2_decap_8
XFILLER_58_801 VPWR VGND sg13g2_fill_1
X_09965_ _04059_ VPWR _01218_ VGND _03995_ _04054_ sg13g2_o21ai_1
X_08916_ _03081_ _03102_ _03103_ VPWR VGND sg13g2_nor2_1
XFILLER_103_268 VPWR VGND sg13g2_decap_8
XFILLER_98_981 VPWR VGND sg13g2_decap_8
XFILLER_69_160 VPWR VGND sg13g2_fill_2
XFILLER_58_812 VPWR VGND sg13g2_fill_1
X_09896_ VPWR _03993_ _03992_ VGND sg13g2_inv_1
X_08847_ _03033_ VPWR _03034_ VGND net1789 _03002_ sg13g2_o21ai_1
XFILLER_100_986 VPWR VGND sg13g2_decap_8
XFILLER_84_163 VPWR VGND sg13g2_fill_1
XFILLER_73_826 VPWR VGND sg13g2_decap_4
XFILLER_72_303 VPWR VGND sg13g2_fill_2
XFILLER_45_506 VPWR VGND sg13g2_decap_8
X_08778_ VPWR _02965_ acc_sub.reg3en.q\[0\] VGND sg13g2_inv_1
XFILLER_27_56 VPWR VGND sg13g2_decap_8
X_07729_ _02035_ _02006_ acc_sub.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_53_561 VPWR VGND sg13g2_decap_8
XFILLER_40_200 VPWR VGND sg13g2_fill_1
XFILLER_14_937 VPWR VGND sg13g2_decap_8
X_10740_ _04748_ _04749_ _04751_ _04752_ _04753_ VPWR VGND sg13g2_nor4_1
XFILLER_80_391 VPWR VGND sg13g2_fill_1
XFILLER_13_436 VPWR VGND sg13g2_fill_1
XFILLER_13_447 VPWR VGND sg13g2_fill_1
X_10671_ _04677_ _04683_ _04674_ _04684_ VPWR VGND sg13g2_nand3_1
X_12410_ _06256_ net1864 _06255_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_77 VPWR VGND sg13g2_decap_8
XFILLER_127_806 VPWR VGND sg13g2_decap_8
X_13390_ VGND VPWR _07006_ net1693 _00806_ _07071_ sg13g2_a21oi_1
X_12341_ _06187_ _06186_ _06176_ VPWR VGND sg13g2_nand2_1
X_12272_ VPWR _06118_ _05964_ VGND sg13g2_inv_1
XFILLER_4_112 VPWR VGND sg13g2_decap_8
XFILLER_107_541 VPWR VGND sg13g2_decap_4
XFILLER_104_0 VPWR VGND sg13g2_fill_2
X_11223_ _05189_ acc_sum.exp_mant_logic0.a\[2\] net1680 acc_sum.op_sign_logic0.mantisa_a\[5\]
+ net1759 VPWR VGND sg13g2_a22oi_1
X_14011_ VPWR _00562_ net21 VGND sg13g2_inv_1
XFILLER_5_679 VPWR VGND sg13g2_fill_1
XFILLER_4_49 VPWR VGND sg13g2_decap_8
X_11154_ net1663 _05123_ _05124_ VPWR VGND sg13g2_nor2b_2
X_11085_ _05060_ _05049_ acc_sum.exp_mant_logic0.b\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_68_96 VPWR VGND sg13g2_fill_1
XFILLER_68_85 VPWR VGND sg13g2_decap_4
XFILLER_68_74 VPWR VGND sg13g2_decap_8
XFILLER_0_351 VPWR VGND sg13g2_decap_8
XFILLER_1_885 VPWR VGND sg13g2_decap_8
X_10105_ _04189_ net1662 _04188_ VPWR VGND sg13g2_nand2_2
XFILLER_103_791 VPWR VGND sg13g2_fill_1
X_14913_ _00714_ VGND VPWR _01433_ acc_sub.seg_reg0.q\[23\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_76_653 VPWR VGND sg13g2_decap_4
XFILLER_48_344 VPWR VGND sg13g2_fill_2
XFILLER_48_333 VPWR VGND sg13g2_decap_8
X_10036_ _04124_ net1662 _04123_ VPWR VGND sg13g2_nand2_2
XFILLER_124_91 VPWR VGND sg13g2_decap_8
XFILLER_91_612 VPWR VGND sg13g2_fill_1
XFILLER_75_141 VPWR VGND sg13g2_fill_2
X_14844_ _00645_ VGND VPWR _01368_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[6\] clknet_leaf_116_clk
+ sg13g2_dfrbpq_2
XFILLER_17_731 VPWR VGND sg13g2_decap_4
X_14775_ _00576_ VGND VPWR _01299_ acc_sub.y\[4\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_11987_ fpmul.reg_b_out\[8\] fpmul.reg_a_out\[8\] _05841_ VPWR VGND sg13g2_xor2_1
XFILLER_17_753 VPWR VGND sg13g2_decap_8
X_13726_ VPWR _00277_ net64 VGND sg13g2_inv_1
X_10938_ _04742_ _04825_ _04945_ VPWR VGND sg13g2_nor2_1
XFILLER_32_734 VPWR VGND sg13g2_decap_8
XFILLER_16_285 VPWR VGND sg13g2_decap_8
XFILLER_31_233 VPWR VGND sg13g2_fill_1
XFILLER_32_745 VPWR VGND sg13g2_fill_1
X_13657_ VPWR _00208_ net68 VGND sg13g2_inv_1
X_10869_ VGND VPWR net1772 _04880_ _04881_ _04771_ sg13g2_a21oi_1
X_12608_ _06424_ fpdiv.div_out\[11\] fpdiv.div_out\[3\] VPWR VGND sg13g2_nand2_1
X_13588_ VPWR _00139_ net124 VGND sg13g2_inv_1
XFILLER_9_941 VPWR VGND sg13g2_decap_8
XFILLER_31_299 VPWR VGND sg13g2_fill_2
XFILLER_118_817 VPWR VGND sg13g2_decap_8
X_12539_ _05378_ _05380_ _05372_ _06356_ VPWR VGND _02722_ sg13g2_nand4_1
XFILLER_8_462 VPWR VGND sg13g2_decap_8
X_14209_ VPWR _00760_ net133 VGND sg13g2_inv_1
XFILLER_99_701 VPWR VGND sg13g2_decap_8
XFILLER_126_883 VPWR VGND sg13g2_decap_8
XFILLER_125_382 VPWR VGND sg13g2_fill_2
XFILLER_98_211 VPWR VGND sg13g2_decap_8
XFILLER_63_1007 VPWR VGND sg13g2_decap_8
XFILLER_99_767 VPWR VGND sg13g2_fill_1
XFILLER_99_756 VPWR VGND sg13g2_decap_8
X_09750_ _03865_ VPWR _03866_ VGND _03832_ _03861_ sg13g2_o21ai_1
XFILLER_98_277 VPWR VGND sg13g2_decap_8
XFILLER_98_266 VPWR VGND sg13g2_fill_1
X_09681_ _03797_ _03796_ net1807 VPWR VGND sg13g2_nand2_1
X_08701_ VGND VPWR net1671 _02841_ _02914_ net1740 sg13g2_a21oi_1
XFILLER_95_995 VPWR VGND sg13g2_decap_8
X_08632_ _02853_ VPWR _02854_ VGND _02746_ _02852_ sg13g2_o21ai_1
XFILLER_55_826 VPWR VGND sg13g2_fill_1
X_08563_ _02786_ VPWR _02787_ VGND _02746_ _02785_ sg13g2_o21ai_1
X_08494_ _02721_ fpdiv.divider0.remainder_reg\[5\] net1708 net1748 fpdiv.divider0.dividend\[5\]
+ VPWR VGND sg13g2_a22oi_1
X_07514_ VPWR VGND _01793_ _01788_ _01835_ _01783_ _01836_ _01791_ sg13g2_a221oi_1
XFILLER_120_49 VPWR VGND sg13g2_decap_8
X_07445_ _01773_ VPWR _01445_ VGND _01772_ net1750 sg13g2_o21ai_1
XFILLER_81_199 VPWR VGND sg13g2_decap_8
Xfanout37 net38 net37 VPWR VGND sg13g2_buf_2
XFILLER_50_520 VPWR VGND sg13g2_decap_8
Xfanout26 net28 net26 VPWR VGND sg13g2_buf_2
XFILLER_22_211 VPWR VGND sg13g2_fill_2
Xfanout15 net72 net15 VPWR VGND sg13g2_buf_2
Xfanout59 net60 net59 VPWR VGND sg13g2_buf_2
Xfanout48 net49 net48 VPWR VGND sg13g2_buf_2
XFILLER_13_14 VPWR VGND sg13g2_decap_8
X_07376_ _01726_ net1886 acc\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_22_288 VPWR VGND sg13g2_decap_8
X_09115_ _03295_ VPWR _03296_ VGND _03167_ _03176_ sg13g2_o21ai_1
XFILLER_109_828 VPWR VGND sg13g2_decap_8
XFILLER_108_305 VPWR VGND sg13g2_fill_1
XFILLER_124_809 VPWR VGND sg13g2_decap_8
X_09046_ net1791 _01715_ _03232_ VPWR VGND sg13g2_nor2_1
XFILLER_123_308 VPWR VGND sg13g2_decap_8
XFILLER_117_872 VPWR VGND sg13g2_decap_8
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_104_533 VPWR VGND sg13g2_decap_4
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_77_439 VPWR VGND sg13g2_fill_1
XFILLER_49_119 VPWR VGND sg13g2_decap_8
X_09948_ _03993_ _04003_ _04044_ VPWR VGND sg13g2_nor2_1
XFILLER_89_299 VPWR VGND sg13g2_decap_4
X_09879_ _03981_ VPWR _01226_ VGND net1768 _03779_ sg13g2_o21ai_1
XFILLER_86_973 VPWR VGND sg13g2_decap_8
XFILLER_73_601 VPWR VGND sg13g2_decap_8
XFILLER_58_675 VPWR VGND sg13g2_decap_8
XFILLER_57_141 VPWR VGND sg13g2_decap_8
XFILLER_46_815 VPWR VGND sg13g2_decap_8
XFILLER_38_77 VPWR VGND sg13g2_decap_8
XFILLER_18_506 VPWR VGND sg13g2_decap_8
XFILLER_18_517 VPWR VGND sg13g2_fill_2
XFILLER_100_794 VPWR VGND sg13g2_decap_8
X_12890_ _06667_ _06666_ fpmul.reg1en.d\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_57_196 VPWR VGND sg13g2_decap_4
X_11910_ net1880 fpmul.seg_reg0.q\[43\] _05784_ VPWR VGND sg13g2_nor2_1
XFILLER_18_539 VPWR VGND sg13g2_fill_1
XFILLER_73_667 VPWR VGND sg13g2_fill_2
XFILLER_54_21 VPWR VGND sg13g2_decap_8
XFILLER_45_358 VPWR VGND sg13g2_decap_4
X_11841_ _05737_ _05739_ _05570_ _05740_ VPWR VGND sg13g2_nand3_1
X_14560_ _00361_ VGND VPWR _01096_ acc_sum.seg_reg0.q\[23\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_61_829 VPWR VGND sg13g2_fill_1
X_11772_ _05676_ _05650_ _05675_ VPWR VGND sg13g2_nand2_1
X_13511_ VPWR _00062_ net37 VGND sg13g2_inv_1
XFILLER_54_98 VPWR VGND sg13g2_fill_1
X_10723_ VPWR _04736_ _04679_ VGND sg13g2_inv_1
X_14491_ _00292_ VGND VPWR net1741 fpdiv.reg2en.q\[0\] clknet_leaf_53_clk sg13g2_dfrbpq_1
X_13442_ _07100_ net1751 sipo.shift_reg\[12\] VPWR VGND sg13g2_nand2_1
X_10654_ VPWR _04667_ _04666_ VGND sg13g2_inv_1
XFILLER_70_86 VPWR VGND sg13g2_fill_2
XFILLER_70_75 VPWR VGND sg13g2_fill_2
X_13373_ _07062_ VPWR _00814_ VGND _06337_ net1694 sg13g2_o21ai_1
X_10585_ _04605_ VPWR _01144_ VGND net1932 _02218_ sg13g2_o21ai_1
XFILLER_10_940 VPWR VGND sg13g2_decap_8
XFILLER_127_636 VPWR VGND sg13g2_decap_8
X_12324_ _06170_ _06160_ _06167_ VPWR VGND sg13g2_xnor2_1
Xclkload29 clknet_leaf_7_clk clkload29/X VPWR VGND sg13g2_buf_8
XFILLER_6_955 VPWR VGND sg13g2_decap_8
Xclkload18 clknet_leaf_144_clk clkload18/X VPWR VGND sg13g2_buf_8
XFILLER_126_168 VPWR VGND sg13g2_decap_8
XFILLER_115_809 VPWR VGND sg13g2_decap_8
XFILLER_5_443 VPWR VGND sg13g2_decap_8
XFILLER_123_820 VPWR VGND sg13g2_decap_8
XFILLER_119_91 VPWR VGND sg13g2_decap_8
XFILLER_114_319 VPWR VGND sg13g2_decap_8
XFILLER_79_62 VPWR VGND sg13g2_decap_8
X_12255_ _06101_ _06098_ _06100_ VPWR VGND sg13g2_nand2_1
XFILLER_79_73 VPWR VGND sg13g2_fill_1
X_11206_ _01090_ _05171_ _05172_ VPWR VGND sg13g2_nand2_1
XFILLER_69_918 VPWR VGND sg13g2_decap_8
X_12186_ _05783_ VPWR _06032_ VGND _05781_ _06031_ sg13g2_o21ai_1
XFILLER_123_897 VPWR VGND sg13g2_decap_8
XFILLER_110_503 VPWR VGND sg13g2_decap_8
XFILLER_1_660 VPWR VGND sg13g2_fill_1
X_11068_ _05045_ VPWR _01101_ VGND _02922_ net1813 sg13g2_o21ai_1
XFILLER_77_962 VPWR VGND sg13g2_decap_8
XFILLER_48_130 VPWR VGND sg13g2_fill_2
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_37_848 VPWR VGND sg13g2_fill_2
X_10019_ _04107_ net1689 _04014_ VPWR VGND sg13g2_nand2_1
X_14827_ _00628_ VGND VPWR _01351_ fpdiv.divider0.remainder_reg\[6\] clknet_leaf_74_clk
+ sg13g2_dfrbpq_2
XFILLER_91_464 VPWR VGND sg13g2_decap_8
XFILLER_91_453 VPWR VGND sg13g2_fill_1
XFILLER_52_818 VPWR VGND sg13g2_decap_8
XFILLER_51_306 VPWR VGND sg13g2_decap_8
XFILLER_17_583 VPWR VGND sg13g2_fill_2
X_14758_ _00559_ VGND VPWR _01282_ acc_sum.exp_mant_logic0.b\[3\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
XFILLER_51_339 VPWR VGND sg13g2_decap_8
X_13709_ VPWR _00260_ net64 VGND sg13g2_inv_1
X_14689_ _00490_ VGND VPWR _01217_ fp16_res_pipe.seg_reg0.q\[26\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
X_07230_ _01600_ VPWR _01601_ VGND _01562_ _01560_ sg13g2_o21ai_1
XFILLER_20_748 VPWR VGND sg13g2_fill_2
X_07161_ VPWR _01533_ acc_sub.op_sign_logic0.mantisa_b\[5\] VGND sg13g2_inv_1
XFILLER_118_625 VPWR VGND sg13g2_fill_2
XFILLER_9_771 VPWR VGND sg13g2_fill_2
XFILLER_8_281 VPWR VGND sg13g2_decap_8
XFILLER_117_168 VPWR VGND sg13g2_decap_8
XFILLER_114_853 VPWR VGND sg13g2_decap_8
XFILLER_113_341 VPWR VGND sg13g2_fill_2
XFILLER_5_70 VPWR VGND sg13g2_decap_8
X_09802_ _03836_ _03859_ _03916_ VPWR VGND sg13g2_nor2_1
XFILLER_87_737 VPWR VGND sg13g2_decap_8
XFILLER_59_428 VPWR VGND sg13g2_decap_4
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
XFILLER_115_49 VPWR VGND sg13g2_decap_8
XFILLER_101_547 VPWR VGND sg13g2_decap_8
X_07994_ fp16_sum_pipe.exp_mant_logic0.a\[4\] _02261_ VPWR VGND sg13g2_inv_4
X_09733_ _03848_ VPWR _03849_ VGND _02928_ _03828_ sg13g2_o21ai_1
X_09664_ _03757_ _03765_ _03780_ _03781_ VPWR VGND sg13g2_nor3_1
XFILLER_83_932 VPWR VGND sg13g2_decap_8
XFILLER_55_612 VPWR VGND sg13g2_fill_2
XFILLER_39_174 VPWR VGND sg13g2_decap_8
XFILLER_39_163 VPWR VGND sg13g2_decap_8
XFILLER_27_325 VPWR VGND sg13g2_decap_8
XFILLER_28_859 VPWR VGND sg13g2_decap_8
X_09595_ _03712_ _02806_ _02918_ acc_sum.add_renorm0.mantisa\[3\] _03670_ VPWR VGND
+ sg13g2_a22oi_1
X_08615_ _02799_ _02837_ _02838_ VPWR VGND sg13g2_nor2_1
XFILLER_82_453 VPWR VGND sg13g2_fill_2
XFILLER_54_144 VPWR VGND sg13g2_decap_8
XFILLER_15_509 VPWR VGND sg13g2_fill_2
XFILLER_27_336 VPWR VGND sg13g2_fill_1
XFILLER_70_637 VPWR VGND sg13g2_decap_4
XFILLER_70_626 VPWR VGND sg13g2_fill_1
XFILLER_42_306 VPWR VGND sg13g2_decap_4
X_08546_ VPWR _02770_ acc_sum.op_sign_logic0.mantisa_b\[4\] VGND sg13g2_inv_1
XFILLER_70_648 VPWR VGND sg13g2_fill_2
XFILLER_42_339 VPWR VGND sg13g2_decap_8
XFILLER_36_892 VPWR VGND sg13g2_decap_8
XFILLER_35_380 VPWR VGND sg13g2_fill_2
X_08477_ _02707_ _02692_ _02706_ VPWR VGND sg13g2_nand2_1
XFILLER_24_35 VPWR VGND sg13g2_decap_8
X_07428_ _01762_ net1749 fpdiv.divider0.divisor\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_50_372 VPWR VGND sg13g2_fill_2
XFILLER_11_726 VPWR VGND sg13g2_decap_8
XFILLER_11_737 VPWR VGND sg13g2_fill_2
X_07359_ _01715_ acc_sub.add_renorm0.exp\[4\] VPWR VGND sg13g2_inv_2
XFILLER_10_236 VPWR VGND sg13g2_fill_2
XFILLER_108_113 VPWR VGND sg13g2_fill_2
XFILLER_108_146 VPWR VGND sg13g2_decap_8
XFILLER_40_56 VPWR VGND sg13g2_decap_8
XFILLER_3_903 VPWR VGND sg13g2_decap_8
X_10370_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[2\] _04419_ _04420_ VPWR VGND sg13g2_nor2_2
XFILLER_124_639 VPWR VGND sg13g2_decap_8
XFILLER_123_105 VPWR VGND sg13g2_decap_8
X_09029_ _03215_ _03192_ _03214_ VPWR VGND sg13g2_nand2_1
XFILLER_2_402 VPWR VGND sg13g2_decap_8
XFILLER_104_341 VPWR VGND sg13g2_decap_8
X_12040_ _05886_ _05884_ _05885_ VPWR VGND sg13g2_nand2_1
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_2_479 VPWR VGND sg13g2_decap_8
XFILLER_120_834 VPWR VGND sg13g2_decap_8
XFILLER_77_247 VPWR VGND sg13g2_fill_1
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_105_60 VPWR VGND sg13g2_decap_8
XFILLER_65_409 VPWR VGND sg13g2_decap_4
X_13991_ VPWR _00542_ net9 VGND sg13g2_inv_1
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_85_280 VPWR VGND sg13g2_fill_2
X_12942_ _06713_ _06714_ _06704_ _00897_ VPWR VGND sg13g2_nand3_1
XFILLER_65_42 VPWR VGND sg13g2_fill_1
XFILLER_19_848 VPWR VGND sg13g2_fill_1
XFILLER_65_64 VPWR VGND sg13g2_decap_4
XFILLER_45_133 VPWR VGND sg13g2_decap_8
X_12873_ acc\[8\] net1908 net1767 _06651_ VPWR VGND sg13g2_nand3_1
X_14612_ _00413_ VGND VPWR _01144_ fp16_sum_pipe.exp_mant_logic0.a\[7\] clknet_leaf_123_clk
+ sg13g2_dfrbpq_2
XFILLER_121_70 VPWR VGND sg13g2_decap_8
XFILLER_26_391 VPWR VGND sg13g2_fill_2
X_11824_ _05724_ _05599_ _05723_ VPWR VGND sg13g2_nand2b_1
XFILLER_81_30 VPWR VGND sg13g2_fill_2
X_14543_ _00344_ VGND VPWR _01079_ acc_sum.op_sign_logic0.mantisa_b\[6\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
XFILLER_42_873 VPWR VGND sg13g2_fill_1
X_11755_ VPWR _05659_ _05658_ VGND sg13g2_inv_1
X_14474_ _00275_ VGND VPWR fpdiv.divider0.en_r fpdiv.divider0.state clknet_leaf_73_clk
+ sg13g2_dfrbpq_2
X_10706_ _04719_ _04681_ _04675_ VPWR VGND sg13g2_nand2b_1
X_13425_ _07091_ VPWR _00791_ VGND _07003_ net1719 sg13g2_o21ai_1
X_11686_ fp16_sum_pipe.add_renorm0.exp\[3\] _05583_ _05590_ VPWR VGND sg13g2_nor2_1
XFILLER_127_433 VPWR VGND sg13g2_decap_8
Xclkload107 clknet_leaf_66_clk clkload107/X VPWR VGND sg13g2_buf_8
X_10637_ fp16_res_pipe.add_renorm0.mantisa\[8\] fp16_res_pipe.add_renorm0.mantisa\[7\]
+ _04646_ _04650_ VPWR VGND sg13g2_nand3_1
XFILLER_10_770 VPWR VGND sg13g2_fill_2
XFILLER_127_444 VPWR VGND sg13g2_decap_8
Xplace1908 load_en net1908 VPWR VGND sg13g2_buf_2
X_13356_ _07052_ net1724 fp16_res_pipe.x2\[2\] VPWR VGND sg13g2_nand2_1
X_10568_ fp16_sum_pipe.exp_mant_logic0.a\[15\] net1931 _04597_ VPWR VGND sg13g2_nor2_1
XFILLER_127_499 VPWR VGND sg13g2_decap_8
XFILLER_114_105 VPWR VGND sg13g2_decap_8
X_13287_ VGND VPWR net1677 _07001_ _00840_ _07002_ sg13g2_a21oi_1
X_12307_ _06062_ _06152_ _06153_ VPWR VGND sg13g2_nor2_1
Xplace1919 net1912 net1919 VPWR VGND sg13g2_buf_2
X_10499_ net1847 fp16_sum_pipe.add_renorm0.mantisa\[7\] _04544_ VPWR VGND sg13g2_nor2_1
X_12238_ _06083_ _06079_ _06084_ VPWR VGND sg13g2_xor2_1
XFILLER_123_661 VPWR VGND sg13g2_fill_2
XFILLER_122_182 VPWR VGND sg13g2_decap_8
XFILLER_111_845 VPWR VGND sg13g2_decap_8
XFILLER_96_534 VPWR VGND sg13g2_decap_8
XFILLER_69_759 VPWR VGND sg13g2_fill_2
X_12169_ _06015_ fpmul.reg_b_out\[2\] VPWR VGND sg13g2_inv_2
XFILLER_96_589 VPWR VGND sg13g2_decap_8
XFILLER_84_729 VPWR VGND sg13g2_decap_8
XFILLER_49_450 VPWR VGND sg13g2_decap_8
XFILLER_65_921 VPWR VGND sg13g2_decap_8
XFILLER_37_612 VPWR VGND sg13g2_fill_2
XFILLER_92_740 VPWR VGND sg13g2_decap_8
XFILLER_37_645 VPWR VGND sg13g2_fill_2
X_08400_ _02636_ VPWR _01359_ VGND _02589_ _02635_ sg13g2_o21ai_1
XFILLER_64_475 VPWR VGND sg13g2_fill_2
XFILLER_36_177 VPWR VGND sg13g2_decap_8
XFILLER_91_294 VPWR VGND sg13g2_fill_1
XFILLER_80_979 VPWR VGND sg13g2_fill_2
XFILLER_80_957 VPWR VGND sg13g2_fill_1
XFILLER_80_946 VPWR VGND sg13g2_decap_8
X_09380_ _03528_ net1674 _03493_ VPWR VGND sg13g2_nand2_1
XFILLER_18_892 VPWR VGND sg13g2_decap_8
XFILLER_24_339 VPWR VGND sg13g2_fill_1
X_08331_ _02576_ _02575_ _02571_ VPWR VGND sg13g2_nand2_2
XFILLER_33_873 VPWR VGND sg13g2_decap_8
XFILLER_60_692 VPWR VGND sg13g2_decap_8
X_08262_ _02510_ _02511_ _02512_ VPWR VGND sg13g2_nor2b_1
XFILLER_119_912 VPWR VGND sg13g2_decap_8
X_07213_ acc_sub.op_sign_logic0.mantisa_b\[0\] acc_sub.op_sign_logic0.mantisa_a\[0\]
+ _01585_ VPWR VGND sg13g2_nor2b_1
XFILLER_118_411 VPWR VGND sg13g2_decap_8
X_08193_ VPWR _02450_ _02408_ VGND sg13g2_inv_1
XFILLER_119_989 VPWR VGND sg13g2_decap_8
X_07144_ VPWR _01516_ _01515_ VGND sg13g2_inv_1
XFILLER_121_609 VPWR VGND sg13g2_decap_8
XFILLER_105_138 VPWR VGND sg13g2_decap_8
XFILLER_105_127 VPWR VGND sg13g2_decap_8
XFILLER_120_119 VPWR VGND sg13g2_decap_8
XFILLER_114_650 VPWR VGND sg13g2_decap_4
XFILLER_113_171 VPWR VGND sg13g2_fill_1
XFILLER_113_160 VPWR VGND sg13g2_decap_8
XFILLER_102_823 VPWR VGND sg13g2_decap_4
XFILLER_102_889 VPWR VGND sg13g2_fill_1
XFILLER_102_878 VPWR VGND sg13g2_decap_8
XFILLER_101_366 VPWR VGND sg13g2_decap_8
XFILLER_59_269 VPWR VGND sg13g2_decap_8
XFILLER_47_409 VPWR VGND sg13g2_decap_8
XFILLER_19_35 VPWR VGND sg13g2_decap_8
X_07977_ _02179_ _02244_ _02250_ VPWR VGND sg13g2_nor2_2
X_09716_ VGND VPWR _03831_ _03832_ _03820_ net1690 sg13g2_a21oi_2
XFILLER_71_902 VPWR VGND sg13g2_decap_8
XFILLER_67_280 VPWR VGND sg13g2_decap_8
XFILLER_28_656 VPWR VGND sg13g2_fill_2
X_09647_ _03764_ _03763_ net1802 VPWR VGND sg13g2_nand2_1
XFILLER_55_475 VPWR VGND sg13g2_decap_8
X_09578_ _03695_ net1806 acc_sum.add_renorm0.mantisa\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_82_283 VPWR VGND sg13g2_fill_2
XFILLER_43_637 VPWR VGND sg13g2_fill_2
XFILLER_35_56 VPWR VGND sg13g2_decap_8
XFILLER_15_328 VPWR VGND sg13g2_decap_4
X_08529_ _02750_ _02752_ _02753_ VPWR VGND sg13g2_nor2_1
XFILLER_70_478 VPWR VGND sg13g2_fill_1
XFILLER_42_147 VPWR VGND sg13g2_decap_4
XFILLER_51_670 VPWR VGND sg13g2_fill_1
XFILLER_11_523 VPWR VGND sg13g2_decap_8
X_11540_ _05445_ _05438_ _05439_ VPWR VGND sg13g2_nand2_1
XFILLER_23_361 VPWR VGND sg13g2_decap_8
XFILLER_23_372 VPWR VGND sg13g2_fill_1
XFILLER_50_180 VPWR VGND sg13g2_fill_1
XFILLER_7_505 VPWR VGND sg13g2_fill_1
XFILLER_109_411 VPWR VGND sg13g2_fill_1
X_11471_ fpdiv.reg_b_out\[10\] fp16_res_pipe.x2\[10\] net1940 _01039_ VPWR VGND sg13g2_mux2_1
XFILLER_51_88 VPWR VGND sg13g2_decap_8
X_14190_ VPWR _00741_ net101 VGND sg13g2_inv_1
X_13210_ _06941_ sipo.word\[0\] VPWR VGND sg13g2_inv_2
X_10422_ _04471_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[7\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[7\]
+ VPWR VGND sg13g2_nand2_1
X_13141_ _06892_ _06891_ _06570_ VPWR VGND sg13g2_nand2b_1
XFILLER_3_700 VPWR VGND sg13g2_fill_1
X_10353_ _04403_ _04402_ VPWR VGND sg13g2_inv_2
X_13072_ _06839_ VPWR _00892_ VGND net1861 _06586_ sg13g2_o21ai_1
X_12023_ net1873 fpmul.seg_reg0.q\[18\] _05872_ VPWR VGND sg13g2_nor2_1
XFILLER_3_777 VPWR VGND sg13g2_fill_2
XFILLER_2_243 VPWR VGND sg13g2_fill_2
XFILLER_2_265 VPWR VGND sg13g2_decap_8
X_10284_ _04298_ _04175_ _04353_ VPWR VGND sg13g2_nor2_1
XFILLER_93_526 VPWR VGND sg13g2_fill_2
XFILLER_93_515 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_fill_2
XFILLER_93_559 VPWR VGND sg13g2_decap_8
XFILLER_46_442 VPWR VGND sg13g2_fill_2
X_13974_ VPWR _00525_ net17 VGND sg13g2_inv_1
XFILLER_74_784 VPWR VGND sg13g2_fill_2
X_12925_ VPWR _06699_ fpmul.reg_p_out\[4\] VGND sg13g2_inv_1
XFILLER_19_678 VPWR VGND sg13g2_decap_8
X_12856_ _06636_ _06635_ net1732 VPWR VGND sg13g2_nand2_1
XFILLER_34_659 VPWR VGND sg13g2_decap_8
XFILLER_18_199 VPWR VGND sg13g2_fill_2
XFILLER_92_84 VPWR VGND sg13g2_decap_4
XFILLER_92_73 VPWR VGND sg13g2_fill_2
XFILLER_61_456 VPWR VGND sg13g2_decap_4
X_11807_ _05708_ _05642_ _05604_ VPWR VGND sg13g2_nand2_1
XFILLER_33_147 VPWR VGND sg13g2_decap_8
X_14526_ _00327_ VGND VPWR _01062_ fpdiv.div_out\[1\] clknet_leaf_72_clk sg13g2_dfrbpq_1
X_11738_ _05634_ _05641_ _05642_ VPWR VGND sg13g2_nor2_2
XFILLER_14_394 VPWR VGND sg13g2_decap_8
X_14457_ _00258_ VGND VPWR _00996_ fpmul.seg_reg0.q\[42\] clknet_leaf_99_clk sg13g2_dfrbpq_1
X_14388_ _00189_ VGND VPWR _00927_ div_result\[1\] clknet_leaf_76_clk sg13g2_dfrbpq_1
X_13408_ _07082_ VPWR _00799_ VGND _07034_ _07076_ sg13g2_o21ai_1
XFILLER_127_252 VPWR VGND sg13g2_decap_8
XFILLER_116_926 VPWR VGND sg13g2_decap_8
Xplace1705 _02654_ net1705 VPWR VGND sg13g2_buf_2
Xplace1716 _06574_ net1716 VPWR VGND sg13g2_buf_1
X_13339_ VPWR _07042_ sipo.word\[9\] VGND sg13g2_inv_1
Xplace1727 _05583_ net1727 VPWR VGND sg13g2_buf_2
XFILLER_6_571 VPWR VGND sg13g2_decap_4
Xplace1749 net1748 net1749 VPWR VGND sg13g2_buf_1
Xplace1738 _03365_ net1738 VPWR VGND sg13g2_buf_2
XFILLER_124_970 VPWR VGND sg13g2_decap_8
X_08880_ _03066_ VPWR _03067_ VGND net1788 _02974_ sg13g2_o21ai_1
XFILLER_97_821 VPWR VGND sg13g2_fill_2
XFILLER_69_534 VPWR VGND sg13g2_fill_2
X_07900_ fp16_sum_pipe.op_sign_logic0.s_a fp16_sum_pipe.exp_mant_logic0.a\[15\] fp16_sum_pipe.reg1en.q\[0\]
+ _01393_ VPWR VGND sg13g2_mux2_1
XFILLER_111_642 VPWR VGND sg13g2_fill_2
X_07831_ _02127_ _02018_ net1747 VPWR VGND sg13g2_nand2_1
XFILLER_110_174 VPWR VGND sg13g2_decap_8
XFILLER_56_228 VPWR VGND sg13g2_fill_2
XFILLER_38_932 VPWR VGND sg13g2_decap_8
X_07762_ _02065_ net1640 _02061_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_431 VPWR VGND sg13g2_decap_8
X_09501_ _03618_ VPWR _01241_ VGND net1916 _03617_ sg13g2_o21ai_1
XFILLER_112_28 VPWR VGND sg13g2_decap_8
X_07693_ _02001_ _01935_ acc_sub.exp_mant_logic0.a\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_64_261 VPWR VGND sg13g2_decap_8
XFILLER_52_401 VPWR VGND sg13g2_decap_8
XFILLER_38_987 VPWR VGND sg13g2_decap_8
XFILLER_37_497 VPWR VGND sg13g2_fill_2
X_09432_ _03573_ VPWR _01265_ VGND fp16_res_pipe.reg2en.q\[0\] _03572_ sg13g2_o21ai_1
XFILLER_25_648 VPWR VGND sg13g2_decap_8
XFILLER_80_787 VPWR VGND sg13g2_fill_2
XFILLER_80_776 VPWR VGND sg13g2_fill_2
XFILLER_40_607 VPWR VGND sg13g2_fill_1
X_09363_ _03513_ net1674 _03496_ VPWR VGND sg13g2_nand2b_1
XFILLER_12_309 VPWR VGND sg13g2_decap_8
X_08314_ _02559_ state\[3\] VPWR VGND sg13g2_inv_2
XFILLER_21_832 VPWR VGND sg13g2_decap_8
X_09294_ fp16_res_pipe.op_sign_logic0.mantisa_b\[0\] fp16_res_pipe.op_sign_logic0.mantisa_a\[0\]
+ _03448_ VPWR VGND sg13g2_nor2b_1
X_08245_ _01368_ _02495_ _02496_ VPWR VGND sg13g2_nand2_1
XFILLER_20_364 VPWR VGND sg13g2_decap_8
X_08176_ _02270_ _02340_ _02434_ VPWR VGND sg13g2_nor2_1
XFILLER_21_14 VPWR VGND sg13g2_decap_8
XFILLER_119_786 VPWR VGND sg13g2_decap_8
XFILLER_118_252 VPWR VGND sg13g2_decap_8
X_07127_ VPWR _01499_ acc_sub.op_sign_logic0.mantisa_a\[10\] VGND sg13g2_inv_1
XFILLER_108_7 VPWR VGND sg13g2_decap_8
XFILLER_106_458 VPWR VGND sg13g2_fill_1
XFILLER_121_417 VPWR VGND sg13g2_decap_4
XFILLER_115_970 VPWR VGND sg13g2_decap_8
XFILLER_106_469 VPWR VGND sg13g2_decap_8
XFILLER_82_1010 VPWR VGND sg13g2_decap_4
XFILLER_47_228 VPWR VGND sg13g2_decap_8
XFILLER_28_420 VPWR VGND sg13g2_decap_8
XFILLER_56_762 VPWR VGND sg13g2_decap_4
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_43_401 VPWR VGND sg13g2_decap_4
X_10971_ _04969_ _04970_ _04968_ _04971_ VPWR VGND sg13g2_nand3_1
XFILLER_28_475 VPWR VGND sg13g2_decap_8
XFILLER_29_976 VPWR VGND sg13g2_decap_8
X_12710_ _06435_ VPWR _06517_ VGND _06427_ _06452_ sg13g2_o21ai_1
XFILLER_71_743 VPWR VGND sg13g2_fill_1
XFILLER_70_220 VPWR VGND sg13g2_decap_8
XFILLER_43_423 VPWR VGND sg13g2_fill_2
XFILLER_43_412 VPWR VGND sg13g2_decap_8
X_13690_ VPWR _00241_ net66 VGND sg13g2_inv_1
X_12641_ _06454_ _06456_ _06453_ _06457_ VPWR VGND sg13g2_nand3_1
XFILLER_71_754 VPWR VGND sg13g2_decap_8
XFILLER_15_147 VPWR VGND sg13g2_fill_1
XFILLER_12_810 VPWR VGND sg13g2_decap_8
XFILLER_12_821 VPWR VGND sg13g2_fill_1
X_12572_ _06388_ _06385_ _06384_ VPWR VGND sg13g2_nand2b_1
XFILLER_62_98 VPWR VGND sg13g2_fill_1
XFILLER_62_87 VPWR VGND sg13g2_decap_8
XFILLER_8_803 VPWR VGND sg13g2_decap_4
XFILLER_11_320 VPWR VGND sg13g2_fill_1
X_14311_ _00112_ VGND VPWR _00004_ sipo.word_ready clknet_leaf_22_clk sg13g2_dfrbpq_2
XFILLER_8_825 VPWR VGND sg13g2_decap_8
XFILLER_12_876 VPWR VGND sg13g2_decap_8
X_11523_ _05428_ _05419_ _05427_ VPWR VGND sg13g2_xnor2_1
X_11454_ _05379_ acc_sub.x2\[3\] net1947 VPWR VGND sg13g2_nand2_1
X_14242_ _00043_ VGND VPWR _00793_ instr\[7\] clknet_leaf_20_clk sg13g2_dfrbpq_1
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_11_397 VPWR VGND sg13g2_decap_4
XFILLER_125_701 VPWR VGND sg13g2_decap_8
X_10405_ _04451_ _04454_ _04455_ VPWR VGND sg13g2_nor2_1
XFILLER_125_767 VPWR VGND sg13g2_decap_8
XFILLER_113_907 VPWR VGND sg13g2_decap_8
X_14173_ VPWR _00724_ net131 VGND sg13g2_inv_1
XFILLER_109_285 VPWR VGND sg13g2_fill_1
X_11385_ _05335_ _05256_ _05334_ VPWR VGND sg13g2_nand2_1
XFILLER_124_266 VPWR VGND sg13g2_decap_8
XFILLER_112_406 VPWR VGND sg13g2_decap_4
X_13124_ _06777_ VPWR _06878_ VGND _06795_ _06799_ sg13g2_o21ai_1
XFILLER_11_91 VPWR VGND sg13g2_decap_8
XFILLER_127_91 VPWR VGND sg13g2_decap_8
XFILLER_106_992 VPWR VGND sg13g2_decap_8
Xclkbuf_4_9_0_clk clknet_0_clk clknet_4_9_0_clk VPWR VGND sg13g2_buf_8
X_13055_ fpmul.seg_reg0.q\[53\] fpmul.seg_reg0.q\[52\] fpmul.seg_reg0.q\[51\] _06823_
+ VPWR VGND sg13g2_nor3_1
XFILLER_3_574 VPWR VGND sg13g2_fill_2
X_10267_ _04336_ VPWR _04337_ VGND _04302_ _04222_ sg13g2_o21ai_1
XFILLER_121_973 VPWR VGND sg13g2_decap_8
X_12006_ net1875 fpmul.seg_reg0.q\[23\] _05860_ VPWR VGND sg13g2_nor2_1
XFILLER_39_707 VPWR VGND sg13g2_fill_2
XFILLER_23_7 VPWR VGND sg13g2_decap_8
XFILLER_93_301 VPWR VGND sg13g2_fill_2
XFILLER_78_375 VPWR VGND sg13g2_fill_2
X_10198_ _04275_ net1829 net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[9\] _03988_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_93_334 VPWR VGND sg13g2_decap_4
XFILLER_47_751 VPWR VGND sg13g2_decap_8
X_13957_ VPWR _00508_ net79 VGND sg13g2_inv_1
XFILLER_81_529 VPWR VGND sg13g2_fill_1
XFILLER_59_1012 VPWR VGND sg13g2_fill_2
XFILLER_19_453 VPWR VGND sg13g2_decap_8
XFILLER_62_743 VPWR VGND sg13g2_fill_2
X_12908_ VGND VPWR net1936 add_result\[5\] _06683_ net1950 sg13g2_a21oi_1
XFILLER_46_283 VPWR VGND sg13g2_fill_1
XFILLER_35_946 VPWR VGND sg13g2_decap_8
XFILLER_34_434 VPWR VGND sg13g2_fill_2
XFILLER_62_765 VPWR VGND sg13g2_fill_1
XFILLER_62_754 VPWR VGND sg13g2_decap_8
XFILLER_61_231 VPWR VGND sg13g2_decap_8
X_13888_ VPWR _00439_ net49 VGND sg13g2_inv_1
X_12839_ _06620_ _06616_ _06619_ _06488_ net1941 VPWR VGND sg13g2_a22oi_1
XFILLER_15_681 VPWR VGND sg13g2_decap_8
X_14509_ _00310_ VGND VPWR _01045_ fpdiv.divider0.dividend\[4\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_1
X_08030_ VGND VPWR net1692 _02282_ _02296_ _02295_ sg13g2_a21oi_1
XFILLER_115_266 VPWR VGND sg13g2_decap_8
XFILLER_104_929 VPWR VGND sg13g2_decap_8
XFILLER_89_629 VPWR VGND sg13g2_decap_8
X_09981_ fp16_res_pipe.exp_mant_logic0.a\[14\] fp16_res_pipe.exp_mant_logic0.a\[13\]
+ fp16_res_pipe.exp_mant_logic0.a\[12\] fp16_res_pipe.exp_mant_logic0.a\[11\] _04070_
+ VPWR VGND sg13g2_nor4_1
X_08932_ _03114_ _03118_ acc_sub.seg_reg1.q\[21\] _03119_ VPWR VGND sg13g2_mux2_1
XFILLER_88_128 VPWR VGND sg13g2_decap_4
X_08863_ _03049_ VPWR _03050_ VGND _02979_ _02997_ sg13g2_o21ai_1
XFILLER_96_172 VPWR VGND sg13g2_fill_2
XFILLER_96_150 VPWR VGND sg13g2_decap_8
XFILLER_69_386 VPWR VGND sg13g2_decap_8
XFILLER_69_364 VPWR VGND sg13g2_fill_2
XFILLER_57_504 VPWR VGND sg13g2_fill_1
X_08794_ _02981_ _02977_ _02974_ VPWR VGND sg13g2_nand2_1
XFILLER_123_49 VPWR VGND sg13g2_decap_8
X_07814_ _02111_ _02006_ net1747 VPWR VGND sg13g2_nand2_1
XFILLER_96_194 VPWR VGND sg13g2_fill_2
XFILLER_85_879 VPWR VGND sg13g2_fill_2
XFILLER_84_323 VPWR VGND sg13g2_fill_2
XFILLER_57_559 VPWR VGND sg13g2_decap_8
X_07745_ _01751_ _02024_ _02050_ VPWR VGND sg13g2_nor2_1
XFILLER_38_784 VPWR VGND sg13g2_decap_4
XFILLER_65_592 VPWR VGND sg13g2_decap_8
XFILLER_16_14 VPWR VGND sg13g2_decap_8
X_07676_ _01986_ acc_sub.exp_mant_logic0.a\[2\] net1672 acc_sub.op_sign_logic0.mantisa_a\[5\]
+ net1780 VPWR VGND sg13g2_a22oi_1
X_09415_ _03558_ VPWR _03559_ VGND _03417_ net1675 sg13g2_o21ai_1
XFILLER_13_607 VPWR VGND sg13g2_decap_8
XFILLER_25_456 VPWR VGND sg13g2_decap_4
XFILLER_26_968 VPWR VGND sg13g2_decap_8
XFILLER_80_595 VPWR VGND sg13g2_decap_8
XFILLER_41_949 VPWR VGND sg13g2_fill_1
X_09346_ _03498_ _03440_ _03452_ VPWR VGND sg13g2_nand2_1
X_09277_ VPWR _03431_ _03430_ VGND sg13g2_inv_1
XFILLER_21_662 VPWR VGND sg13g2_fill_1
XFILLER_21_673 VPWR VGND sg13g2_decap_8
XFILLER_32_35 VPWR VGND sg13g2_decap_8
X_08228_ _02480_ _02481_ _02479_ _02482_ VPWR VGND sg13g2_nand3_1
XFILLER_107_745 VPWR VGND sg13g2_decap_8
X_08159_ _02419_ fp16_sum_pipe.exp_mant_logic0.a\[0\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[3\]
+ net1776 VPWR VGND sg13g2_a22oi_1
X_11170_ _05139_ _05110_ _05023_ VPWR VGND sg13g2_nand2b_1
XFILLER_121_203 VPWR VGND sg13g2_decap_8
XFILLER_79_128 VPWR VGND sg13g2_decap_8
X_10121_ _04201_ _04202_ _04203_ _04204_ VPWR VGND sg13g2_nor3_1
XFILLER_0_533 VPWR VGND sg13g2_decap_8
X_10052_ _04121_ _04139_ _04105_ _04140_ VPWR VGND sg13g2_nand3_1
XFILLER_103_995 VPWR VGND sg13g2_decap_8
XFILLER_94_109 VPWR VGND sg13g2_fill_1
XFILLER_76_824 VPWR VGND sg13g2_fill_2
XFILLER_0_577 VPWR VGND sg13g2_decap_8
XFILLER_48_537 VPWR VGND sg13g2_decap_8
X_14860_ _00661_ VGND VPWR _01384_ fp16_sum_pipe.seg_reg0.q\[22\] clknet_leaf_121_clk
+ sg13g2_dfrbpq_1
X_13811_ VPWR _00362_ net77 VGND sg13g2_inv_1
XFILLER_75_367 VPWR VGND sg13g2_decap_8
X_14791_ _00592_ VGND VPWR _01315_ acc_sum.exp_mant_logic0.a\[4\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_13742_ VPWR _00293_ net137 VGND sg13g2_inv_1
XFILLER_56_581 VPWR VGND sg13g2_decap_8
XFILLER_44_765 VPWR VGND sg13g2_fill_1
XFILLER_17_968 VPWR VGND sg13g2_decap_8
X_10954_ _04954_ _04952_ _04959_ _04960_ VPWR VGND sg13g2_a21o_1
XFILLER_28_294 VPWR VGND sg13g2_fill_2
X_13673_ VPWR _00224_ net125 VGND sg13g2_inv_1
XFILLER_73_75 VPWR VGND sg13g2_fill_2
XFILLER_71_573 VPWR VGND sg13g2_decap_8
XFILLER_43_275 VPWR VGND sg13g2_decap_8
X_10885_ _04896_ _04892_ _04895_ VPWR VGND sg13g2_nand2_1
X_12624_ _06439_ VPWR _06440_ VGND net1852 fpdiv.div_out\[6\] sg13g2_o21ai_1
XFILLER_12_640 VPWR VGND sg13g2_fill_2
X_12555_ VPWR _06371_ div_result\[14\] VGND sg13g2_inv_1
XFILLER_12_651 VPWR VGND sg13g2_decap_8
X_11506_ _05410_ VPWR _05411_ VGND net1840 _05409_ sg13g2_o21ai_1
XFILLER_12_695 VPWR VGND sg13g2_decap_8
X_12486_ net1872 fpmul.seg_reg0.q\[7\] _06324_ VPWR VGND sg13g2_nor2_1
XFILLER_8_677 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
X_11437_ net1937 fpdiv.reg_a_out\[9\] _05368_ VPWR VGND sg13g2_nor2_1
X_14225_ _00026_ VGND VPWR _00776_ sipo.shift_reg\[6\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_7_198 VPWR VGND sg13g2_fill_2
XFILLER_7_187 VPWR VGND sg13g2_fill_2
X_14156_ VPWR _00707_ net130 VGND sg13g2_inv_1
X_11368_ _05319_ _05211_ net1812 VPWR VGND sg13g2_nand2_1
X_13107_ _06788_ _06774_ _06865_ VPWR VGND sg13g2_xor2_1
XFILLER_3_371 VPWR VGND sg13g2_decap_8
X_10319_ _04377_ net1920 fp16_res_pipe.x2\[6\] VPWR VGND sg13g2_nand2_1
X_14087_ VPWR _00638_ net89 VGND sg13g2_inv_1
X_11299_ _05258_ net1634 _05255_ VPWR VGND sg13g2_nand2b_1
XFILLER_121_770 VPWR VGND sg13g2_decap_8
XFILLER_94_621 VPWR VGND sg13g2_decap_8
XFILLER_78_161 VPWR VGND sg13g2_decap_8
X_13038_ _05873_ _06805_ _06806_ VPWR VGND sg13g2_nor2_1
XFILLER_120_280 VPWR VGND sg13g2_decap_8
XFILLER_78_172 VPWR VGND sg13g2_fill_2
XFILLER_94_665 VPWR VGND sg13g2_decap_8
XFILLER_82_827 VPWR VGND sg13g2_decap_8
XFILLER_82_805 VPWR VGND sg13g2_decap_8
XFILLER_66_356 VPWR VGND sg13g2_decap_8
X_07530_ _01851_ net1782 acc_sub.seg_reg0.q\[27\] VPWR VGND sg13g2_nand2_1
XFILLER_93_186 VPWR VGND sg13g2_decap_8
XFILLER_82_849 VPWR VGND sg13g2_decap_8
XFILLER_81_315 VPWR VGND sg13g2_fill_1
XFILLER_35_721 VPWR VGND sg13g2_decap_8
XFILLER_90_860 VPWR VGND sg13g2_fill_2
XFILLER_23_905 VPWR VGND sg13g2_decap_8
X_07461_ VPWR _01784_ acc_sub.exp_mant_logic0.b\[13\] VGND sg13g2_inv_1
XFILLER_22_426 VPWR VGND sg13g2_fill_2
XFILLER_97_0 VPWR VGND sg13g2_decap_8
X_07392_ _01736_ VPWR _01461_ VGND net1895 _01735_ sg13g2_o21ai_1
X_09200_ _03356_ VPWR _01280_ VGND net1902 _03355_ sg13g2_o21ai_1
XFILLER_34_286 VPWR VGND sg13g2_fill_1
X_09131_ _03311_ _03164_ _03165_ VPWR VGND sg13g2_nand2b_1
X_09062_ _03089_ VPWR _03247_ VGND _03190_ _03246_ sg13g2_o21ai_1
XFILLER_108_509 VPWR VGND sg13g2_decap_8
XFILLER_8_70 VPWR VGND sg13g2_decap_8
X_08013_ VPWR _02279_ _02278_ VGND sg13g2_inv_1
XFILLER_118_49 VPWR VGND sg13g2_decap_8
XFILLER_116_542 VPWR VGND sg13g2_decap_8
XFILLER_104_715 VPWR VGND sg13g2_decap_8
XFILLER_103_214 VPWR VGND sg13g2_fill_1
XFILLER_103_203 VPWR VGND sg13g2_decap_8
XFILLER_98_960 VPWR VGND sg13g2_decap_8
X_09964_ _04059_ fp16_res_pipe.exp_mant_logic0.a\[12\] net1682 net1766 fp16_res_pipe.seg_reg0.q\[27\]
+ VPWR VGND sg13g2_a22oi_1
X_08915_ VGND VPWR _03091_ _03101_ _03102_ net1785 sg13g2_a21oi_1
X_09895_ _03992_ fp16_res_pipe.exp_mant_logic0.a\[14\] fp16_res_pipe.exp_mant_logic0.b\[14\]
+ VPWR VGND sg13g2_xnor2_1
X_08846_ _03033_ net1789 acc_sub.add_renorm0.mantisa\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_69_172 VPWR VGND sg13g2_decap_8
XFILLER_57_334 VPWR VGND sg13g2_decap_4
XFILLER_100_965 VPWR VGND sg13g2_decap_8
XFILLER_84_153 VPWR VGND sg13g2_decap_4
XFILLER_84_142 VPWR VGND sg13g2_fill_1
XFILLER_73_805 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_8
X_08777_ _02964_ VPWR _01311_ VGND net1899 _02963_ sg13g2_o21ai_1
XFILLER_57_389 VPWR VGND sg13g2_decap_8
X_07728_ _02034_ _02018_ acc_sub.exp_mant_logic0.a\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_72_359 VPWR VGND sg13g2_decap_8
XFILLER_53_540 VPWR VGND sg13g2_decap_8
X_07659_ _01968_ _01969_ _01967_ _01970_ VPWR VGND sg13g2_nand3_1
XFILLER_81_882 VPWR VGND sg13g2_fill_2
XFILLER_41_724 VPWR VGND sg13g2_decap_8
XFILLER_14_916 VPWR VGND sg13g2_decap_8
XFILLER_43_56 VPWR VGND sg13g2_decap_8
XFILLER_40_212 VPWR VGND sg13g2_decap_8
XFILLER_9_408 VPWR VGND sg13g2_fill_1
X_10670_ _04683_ _04679_ _04681_ VPWR VGND sg13g2_nand2_1
X_09329_ _03482_ _03361_ net1823 VPWR VGND sg13g2_nand2_1
XFILLER_22_982 VPWR VGND sg13g2_decap_8
X_12340_ _06186_ _06174_ _06179_ VPWR VGND sg13g2_nand2_1
XFILLER_5_614 VPWR VGND sg13g2_decap_8
XFILLER_119_391 VPWR VGND sg13g2_decap_8
X_12271_ VPWR _06117_ _06116_ VGND sg13g2_inv_1
X_11222_ _05188_ _05151_ _05187_ VPWR VGND sg13g2_nand2_1
X_14010_ VPWR _00561_ net19 VGND sg13g2_inv_1
XFILLER_68_20 VPWR VGND sg13g2_fill_2
XFILLER_4_168 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_122_534 VPWR VGND sg13g2_fill_2
X_11153_ _05112_ _05122_ _05123_ VPWR VGND sg13g2_nor2_1
XFILLER_0_330 VPWR VGND sg13g2_decap_8
XFILLER_122_578 VPWR VGND sg13g2_fill_2
XFILLER_89_993 VPWR VGND sg13g2_decap_8
XFILLER_88_470 VPWR VGND sg13g2_decap_4
X_11084_ _05058_ _05059_ _05057_ _01099_ VPWR VGND sg13g2_nand3_1
XFILLER_49_813 VPWR VGND sg13g2_fill_2
XFILLER_1_864 VPWR VGND sg13g2_decap_8
X_10104_ _04111_ _04145_ _04188_ VPWR VGND sg13g2_nor2_1
X_14912_ _00713_ VGND VPWR _01432_ acc_sub.seg_reg0.q\[22\] clknet_leaf_44_clk sg13g2_dfrbpq_1
XFILLER_88_492 VPWR VGND sg13g2_decap_8
XFILLER_76_632 VPWR VGND sg13g2_decap_8
XFILLER_75_120 VPWR VGND sg13g2_decap_8
X_10035_ _04111_ _04122_ _04123_ VPWR VGND sg13g2_nor2_1
XFILLER_124_70 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_48_356 VPWR VGND sg13g2_decap_4
X_14843_ _00644_ VGND VPWR _01367_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[5\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
XFILLER_48_389 VPWR VGND sg13g2_fill_1
XFILLER_1_1013 VPWR VGND sg13g2_fill_1
X_14774_ _00575_ VGND VPWR _01298_ acc_sub.y\[3\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_90_134 VPWR VGND sg13g2_fill_2
X_11986_ fpmul.reg_a_out\[7\] fpmul.reg_b_out\[7\] _05840_ VPWR VGND sg13g2_nor2_1
XFILLER_90_178 VPWR VGND sg13g2_decap_8
XFILLER_71_370 VPWR VGND sg13g2_decap_4
X_13725_ VPWR _00276_ net63 VGND sg13g2_inv_1
X_10937_ VGND VPWR _04694_ _04809_ _04944_ _04943_ sg13g2_a21oi_1
X_13656_ VPWR _00207_ net68 VGND sg13g2_inv_1
X_12607_ _06422_ VPWR _06423_ VGND _06421_ fpdiv.div_out\[4\] sg13g2_o21ai_1
X_10868_ _04880_ _04858_ _04879_ VPWR VGND sg13g2_xnor2_1
XFILLER_9_920 VPWR VGND sg13g2_decap_8
XFILLER_32_779 VPWR VGND sg13g2_decap_4
X_13587_ VPWR _00138_ net121 VGND sg13g2_inv_1
XFILLER_13_982 VPWR VGND sg13g2_decap_8
X_10799_ _04802_ _04810_ _04811_ VPWR VGND sg13g2_nor2_1
X_12538_ _06355_ _05374_ _05376_ VPWR VGND sg13g2_nand2_1
XFILLER_9_997 VPWR VGND sg13g2_decap_8
X_12469_ _06020_ _06057_ _06308_ _06311_ VPWR VGND sg13g2_nand3_1
XFILLER_126_862 VPWR VGND sg13g2_decap_8
X_14208_ VPWR _00759_ net132 VGND sg13g2_inv_1
X_14139_ VPWR _00690_ net89 VGND sg13g2_inv_1
XFILLER_100_206 VPWR VGND sg13g2_fill_2
X_09680_ _03796_ acc_sum.add_renorm0.exp\[5\] _03790_ VPWR VGND sg13g2_xnor2_1
X_08700_ _02913_ net1668 _02842_ VPWR VGND sg13g2_nand2_1
XFILLER_79_481 VPWR VGND sg13g2_decap_8
XFILLER_39_334 VPWR VGND sg13g2_decap_8
XFILLER_95_974 VPWR VGND sg13g2_decap_8
X_08631_ VGND VPWR _02737_ _02740_ _02853_ _02736_ sg13g2_a21oi_1
XFILLER_67_676 VPWR VGND sg13g2_fill_1
XFILLER_66_153 VPWR VGND sg13g2_fill_1
XFILLER_66_131 VPWR VGND sg13g2_decap_8
XFILLER_12_0 VPWR VGND sg13g2_decap_8
XFILLER_81_112 VPWR VGND sg13g2_fill_1
XFILLER_67_687 VPWR VGND sg13g2_fill_2
XFILLER_54_326 VPWR VGND sg13g2_decap_4
X_08562_ VGND VPWR _02737_ _02742_ _02786_ _02735_ sg13g2_a21oi_1
XFILLER_82_657 VPWR VGND sg13g2_fill_1
XFILLER_81_145 VPWR VGND sg13g2_fill_2
XFILLER_70_808 VPWR VGND sg13g2_decap_4
XFILLER_54_359 VPWR VGND sg13g2_decap_8
XFILLER_120_28 VPWR VGND sg13g2_decap_8
X_08493_ _02719_ fpdiv.divider0.remainder_reg\[4\] _02720_ VPWR VGND sg13g2_xor2_1
X_07513_ _01798_ _01834_ _01794_ _01835_ VPWR VGND sg13g2_a21o_1
XFILLER_63_882 VPWR VGND sg13g2_decap_8
X_07444_ _01773_ net1750 fpdiv.divider0.divisor\[5\] VPWR VGND sg13g2_nand2_1
Xfanout38 net39 net38 VPWR VGND sg13g2_buf_2
Xfanout27 net28 net27 VPWR VGND sg13g2_buf_1
Xfanout16 net17 net16 VPWR VGND sg13g2_buf_2
Xfanout49 net72 net49 VPWR VGND sg13g2_buf_1
XFILLER_22_267 VPWR VGND sg13g2_decap_8
XFILLER_109_807 VPWR VGND sg13g2_decap_8
X_07375_ VPWR _01725_ acc_sub.exp_mant_logic0.a\[14\] VGND sg13g2_inv_1
X_09114_ VGND VPWR _03167_ _03176_ _03295_ _03091_ sg13g2_a21oi_1
X_09045_ _03220_ _03230_ _03231_ VPWR VGND sg13g2_nor2_1
XFILLER_108_339 VPWR VGND sg13g2_decap_8
XFILLER_89_19 VPWR VGND sg13g2_fill_1
XFILLER_117_851 VPWR VGND sg13g2_decap_8
XFILLER_116_383 VPWR VGND sg13g2_fill_1
XFILLER_104_523 VPWR VGND sg13g2_decap_4
XFILLER_2_639 VPWR VGND sg13g2_fill_2
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_104_556 VPWR VGND sg13g2_decap_8
XFILLER_77_407 VPWR VGND sg13g2_fill_2
X_09947_ _04042_ VPWR _04043_ VGND _03996_ _04041_ sg13g2_o21ai_1
XFILLER_86_952 VPWR VGND sg13g2_decap_8
X_09878_ _03981_ net1768 acc_sum.y\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_38_56 VPWR VGND sg13g2_decap_8
X_08829_ net1704 _02990_ _02995_ _03016_ VPWR VGND sg13g2_nand3_1
XFILLER_73_635 VPWR VGND sg13g2_decap_8
XFILLER_73_624 VPWR VGND sg13g2_decap_8
XFILLER_72_101 VPWR VGND sg13g2_fill_2
XFILLER_57_175 VPWR VGND sg13g2_fill_1
XFILLER_45_315 VPWR VGND sg13g2_decap_4
XFILLER_72_145 VPWR VGND sg13g2_decap_8
XFILLER_45_337 VPWR VGND sg13g2_decap_8
X_11840_ net1758 VPWR _05739_ VGND _05667_ _05738_ sg13g2_o21ai_1
X_11771_ VGND VPWR net1758 _05674_ _05675_ _05572_ sg13g2_a21oi_1
X_13510_ VPWR _00061_ net84 VGND sg13g2_inv_1
XFILLER_41_521 VPWR VGND sg13g2_decap_8
XFILLER_13_201 VPWR VGND sg13g2_decap_8
X_10722_ VGND VPWR _04720_ _04735_ _04734_ _04722_ sg13g2_a21oi_2
X_14490_ _00291_ VGND VPWR _01028_ add_result\[15\] clknet_leaf_121_clk sg13g2_dfrbpq_2
XFILLER_13_267 VPWR VGND sg13g2_fill_1
X_13441_ _07099_ VPWR _00783_ VGND _06914_ net1751 sg13g2_o21ai_1
X_10653_ _04649_ _04665_ _04666_ VPWR VGND sg13g2_nor2_2
XFILLER_127_604 VPWR VGND sg13g2_decap_8
XFILLER_103_1013 VPWR VGND sg13g2_fill_1
XFILLER_103_1002 VPWR VGND sg13g2_decap_8
X_13372_ _07062_ net1695 sipo.word\[12\] VPWR VGND sg13g2_nand2_1
X_10584_ _04605_ acc_sub.x2\[7\] net1931 VPWR VGND sg13g2_nand2_1
XFILLER_86_1008 VPWR VGND sg13g2_decap_4
X_12323_ _06169_ _06168_ _06159_ VPWR VGND sg13g2_nand2b_1
XFILLER_6_934 VPWR VGND sg13g2_decap_8
XFILLER_5_422 VPWR VGND sg13g2_decap_8
XFILLER_5_400 VPWR VGND sg13g2_decap_8
XFILLER_10_996 VPWR VGND sg13g2_decap_8
Xclkload19 clkload19/Y clknet_leaf_0_clk VPWR VGND sg13g2_inv_2
XFILLER_126_147 VPWR VGND sg13g2_decap_8
XFILLER_119_70 VPWR VGND sg13g2_decap_8
XFILLER_79_30 VPWR VGND sg13g2_fill_2
XFILLER_108_895 VPWR VGND sg13g2_decap_4
X_12254_ VPWR _06100_ _06099_ VGND sg13g2_inv_1
XFILLER_5_499 VPWR VGND sg13g2_decap_8
X_11205_ _05172_ acc_sum.exp_mant_logic0.a\[3\] net1680 acc_sum.op_sign_logic0.mantisa_a\[6\]
+ net1759 VPWR VGND sg13g2_a22oi_1
X_12185_ VPWR _06031_ fpmul.reg_b_out\[6\] VGND sg13g2_inv_1
XFILLER_123_876 VPWR VGND sg13g2_decap_8
XFILLER_96_716 VPWR VGND sg13g2_decap_4
X_11136_ _05106_ _05095_ _05105_ VPWR VGND sg13g2_nand2_2
XFILLER_68_407 VPWR VGND sg13g2_fill_1
XFILLER_77_941 VPWR VGND sg13g2_decap_8
XFILLER_23_1003 VPWR VGND sg13g2_decap_8
XFILLER_95_84 VPWR VGND sg13g2_decap_8
XFILLER_92_900 VPWR VGND sg13g2_fill_2
XFILLER_76_462 VPWR VGND sg13g2_fill_2
X_11067_ _05044_ VPWR _05045_ VGND acc_sum.exp_mant_logic0.b\[13\] _05042_ sg13g2_o21ai_1
XFILLER_37_816 VPWR VGND sg13g2_fill_1
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_91_410 VPWR VGND sg13g2_decap_4
XFILLER_64_635 VPWR VGND sg13g2_decap_8
X_14826_ _00627_ VGND VPWR _01350_ fpdiv.divider0.remainder_reg\[5\] clknet_leaf_74_clk
+ sg13g2_dfrbpq_2
XFILLER_92_988 VPWR VGND sg13g2_decap_8
X_14757_ _00558_ VGND VPWR _01281_ acc_sum.exp_mant_logic0.b\[2\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
X_13708_ VPWR _00259_ net63 VGND sg13g2_inv_1
X_11969_ _05823_ fpmul.reg_a_out\[13\] fpmul.reg_b_out\[13\] VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_137_clk clknet_5_2__leaf_clk clknet_leaf_137_clk VPWR VGND sg13g2_buf_8
XFILLER_60_874 VPWR VGND sg13g2_decap_4
X_14688_ _00489_ VGND VPWR _01216_ fp16_res_pipe.seg_reg0.q\[25\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_1
X_13639_ VPWR _00190_ net124 VGND sg13g2_inv_1
XFILLER_32_598 VPWR VGND sg13g2_decap_8
X_07160_ acc_sub.op_sign_logic0.mantisa_b\[5\] _01531_ _01532_ VPWR VGND sg13g2_nor2_1
XFILLER_118_604 VPWR VGND sg13g2_decap_8
XFILLER_13_790 VPWR VGND sg13g2_fill_1
XFILLER_8_260 VPWR VGND sg13g2_fill_2
XFILLER_9_783 VPWR VGND sg13g2_decap_8
XFILLER_118_659 VPWR VGND sg13g2_fill_2
XFILLER_117_147 VPWR VGND sg13g2_decap_8
XFILLER_126_692 VPWR VGND sg13g2_fill_2
XFILLER_114_832 VPWR VGND sg13g2_decap_8
XFILLER_115_28 VPWR VGND sg13g2_decap_8
XFILLER_113_364 VPWR VGND sg13g2_decap_8
X_09801_ net1803 _03914_ _03912_ _03915_ VPWR VGND sg13g2_nand3_1
XFILLER_101_515 VPWR VGND sg13g2_decap_8
XFILLER_99_587 VPWR VGND sg13g2_decap_4
XFILLER_86_204 VPWR VGND sg13g2_fill_2
XFILLER_101_526 VPWR VGND sg13g2_fill_2
X_09732_ _03848_ _03828_ _03801_ VPWR VGND sg13g2_nand2_1
X_07993_ _02260_ fp16_sum_pipe.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_inv_2
XFILLER_83_911 VPWR VGND sg13g2_decap_8
XFILLER_28_816 VPWR VGND sg13g2_fill_1
X_09663_ _03780_ _03775_ _03779_ VPWR VGND sg13g2_nand2_1
XFILLER_27_304 VPWR VGND sg13g2_decap_8
X_09594_ _03703_ _03710_ _03711_ VPWR VGND sg13g2_nor2_1
X_08614_ _02837_ _02788_ _02836_ _02810_ net1740 VPWR VGND sg13g2_a22oi_1
XFILLER_82_443 VPWR VGND sg13g2_fill_2
XFILLER_43_808 VPWR VGND sg13g2_fill_1
X_08545_ VPWR _02769_ _02768_ VGND sg13g2_inv_1
XFILLER_83_988 VPWR VGND sg13g2_decap_8
XFILLER_42_318 VPWR VGND sg13g2_decap_8
XFILLER_126_1002 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_128_clk clknet_5_6__leaf_clk clknet_leaf_128_clk VPWR VGND sg13g2_buf_8
XFILLER_35_392 VPWR VGND sg13g2_fill_1
XFILLER_24_14 VPWR VGND sg13g2_decap_8
XFILLER_126_1013 VPWR VGND sg13g2_fill_1
X_08476_ _02706_ _02669_ _02668_ VPWR VGND sg13g2_xnor2_1
XFILLER_10_215 VPWR VGND sg13g2_decap_8
X_07358_ _01714_ VPWR _01473_ VGND net1799 _01713_ sg13g2_o21ai_1
XFILLER_40_35 VPWR VGND sg13g2_decap_8
X_07289_ _01656_ _01636_ VPWR VGND sg13g2_inv_2
X_09028_ net1785 _03201_ _03213_ _03214_ VPWR VGND sg13g2_nor3_1
XFILLER_116_180 VPWR VGND sg13g2_decap_8
XFILLER_3_959 VPWR VGND sg13g2_decap_8
XFILLER_120_813 VPWR VGND sg13g2_decap_8
XFILLER_77_204 VPWR VGND sg13g2_fill_1
XFILLER_2_458 VPWR VGND sg13g2_decap_8
XFILLER_78_738 VPWR VGND sg13g2_fill_2
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_59_974 VPWR VGND sg13g2_fill_1
XFILLER_59_963 VPWR VGND sg13g2_decap_8
X_13990_ VPWR _00541_ net9 VGND sg13g2_inv_1
XFILLER_100_581 VPWR VGND sg13g2_decap_8
XFILLER_86_793 VPWR VGND sg13g2_decap_8
X_12941_ _06714_ net1717 _00008_ VPWR VGND sg13g2_nand2_1
X_12872_ VGND VPWR net1935 add_result\[8\] _06650_ net1949 sg13g2_a21oi_1
XFILLER_46_657 VPWR VGND sg13g2_fill_2
XFILLER_46_646 VPWR VGND sg13g2_decap_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
X_14611_ _00412_ VGND VPWR _01143_ fp16_sum_pipe.exp_mant_logic0.a\[6\] clknet_leaf_118_clk
+ sg13g2_dfrbpq_2
XFILLER_27_860 VPWR VGND sg13g2_decap_8
X_11823_ VGND VPWR _05598_ _05444_ _05723_ _05592_ sg13g2_a21oi_1
XFILLER_45_189 VPWR VGND sg13g2_decap_8
XFILLER_26_381 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_119_clk clknet_5_10__leaf_clk clknet_leaf_119_clk VPWR VGND sg13g2_buf_8
X_14542_ _00343_ VGND VPWR _01078_ acc_sum.op_sign_logic0.mantisa_b\[5\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_53_1007 VPWR VGND sg13g2_decap_8
XFILLER_14_554 VPWR VGND sg13g2_decap_8
X_11754_ _05657_ VPWR _05658_ VGND _04465_ _05589_ sg13g2_o21ai_1
X_14473_ _00274_ VGND VPWR _01012_ fpdiv.divider0.counter\[3\] clknet_leaf_72_clk
+ sg13g2_dfrbpq_1
XFILLER_41_384 VPWR VGND sg13g2_fill_2
X_10705_ _04715_ _04712_ _04717_ _04718_ VPWR VGND sg13g2_a21o_1
X_11685_ _05589_ _04589_ _05576_ VPWR VGND sg13g2_xnor2_1
X_13424_ _07091_ net1719 instr\[5\] VPWR VGND sg13g2_nand2_1
X_10636_ VPWR _04649_ _04647_ VGND sg13g2_inv_1
Xclkload108 clknet_leaf_59_clk clkload108/X VPWR VGND sg13g2_buf_8
XFILLER_14_91 VPWR VGND sg13g2_fill_1
X_13355_ _07051_ VPWR _00821_ VGND _07010_ net1723 sg13g2_o21ai_1
Xplace1909 fp16_res_pipe.reg1en.d\[0\] net1909 VPWR VGND sg13g2_buf_2
X_10567_ _04596_ VPWR _01153_ VGND net1844 _04595_ sg13g2_o21ai_1
XFILLER_127_478 VPWR VGND sg13g2_decap_8
X_13286_ acc\[6\] net1677 _07002_ VPWR VGND sg13g2_nor2_1
X_12306_ _06152_ _06149_ _06151_ VPWR VGND sg13g2_nand2_1
XFILLER_53_7 VPWR VGND sg13g2_decap_8
X_10498_ _04543_ _04403_ _04542_ VPWR VGND sg13g2_xnor2_1
XFILLER_107_191 VPWR VGND sg13g2_decap_8
X_12237_ _06081_ _06082_ _06083_ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_14__f_clk clknet_4_7_0_clk clknet_5_14__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_122_161 VPWR VGND sg13g2_decap_8
XFILLER_111_824 VPWR VGND sg13g2_decap_8
XFILLER_110_323 VPWR VGND sg13g2_decap_8
X_12168_ _06014_ _06011_ _06013_ VPWR VGND sg13g2_nand2_1
XFILLER_110_345 VPWR VGND sg13g2_fill_2
XFILLER_84_708 VPWR VGND sg13g2_decap_8
XFILLER_77_760 VPWR VGND sg13g2_fill_1
X_11119_ VGND VPWR _05034_ _05005_ _05089_ _05003_ sg13g2_a21oi_1
X_12099_ _05945_ _05943_ _05944_ VPWR VGND sg13g2_nand2_1
XFILLER_83_229 VPWR VGND sg13g2_fill_1
XFILLER_83_218 VPWR VGND sg13g2_decap_8
XFILLER_77_771 VPWR VGND sg13g2_decap_4
XFILLER_76_281 VPWR VGND sg13g2_decap_8
XFILLER_65_966 VPWR VGND sg13g2_decap_4
XFILLER_36_112 VPWR VGND sg13g2_decap_8
XFILLER_25_808 VPWR VGND sg13g2_fill_2
XFILLER_92_774 VPWR VGND sg13g2_decap_8
XFILLER_52_616 VPWR VGND sg13g2_decap_8
XFILLER_36_156 VPWR VGND sg13g2_decap_8
XFILLER_18_871 VPWR VGND sg13g2_decap_8
X_14809_ _00610_ VGND VPWR _01333_ acc_sum.add_renorm0.exp\[6\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_2
XFILLER_51_137 VPWR VGND sg13g2_decap_4
X_08330_ VPWR _02575_ _02568_ VGND sg13g2_inv_1
XFILLER_60_671 VPWR VGND sg13g2_decap_8
XFILLER_33_885 VPWR VGND sg13g2_fill_1
X_08261_ _02511_ _02347_ net1842 VPWR VGND sg13g2_nand2_1
X_07212_ VPWR _01584_ _01583_ VGND sg13g2_inv_1
XFILLER_32_395 VPWR VGND sg13g2_decap_4
X_08192_ _02269_ _02380_ _02449_ VPWR VGND sg13g2_nor2_1
XFILLER_20_568 VPWR VGND sg13g2_fill_1
XFILLER_119_968 VPWR VGND sg13g2_decap_8
X_07143_ _01508_ _01514_ _01515_ VPWR VGND sg13g2_nor2_1
XFILLER_118_478 VPWR VGND sg13g2_decap_8
XFILLER_106_629 VPWR VGND sg13g2_fill_1
XFILLER_106_618 VPWR VGND sg13g2_decap_8
XFILLER_10_49 VPWR VGND sg13g2_decap_8
XFILLER_126_49 VPWR VGND sg13g2_decap_8
XFILLER_102_813 VPWR VGND sg13g2_decap_4
XFILLER_114_695 VPWR VGND sg13g2_decap_8
XFILLER_113_183 VPWR VGND sg13g2_fill_1
XFILLER_87_513 VPWR VGND sg13g2_fill_2
XFILLER_59_237 VPWR VGND sg13g2_decap_8
XFILLER_101_345 VPWR VGND sg13g2_decap_8
XFILLER_19_14 VPWR VGND sg13g2_decap_8
X_09715_ acc_sum.add_renorm0.exp\[6\] net1690 _03831_ VPWR VGND sg13g2_nor2_1
XFILLER_28_613 VPWR VGND sg13g2_decap_8
X_09646_ _03761_ _03762_ _03760_ _03763_ VPWR VGND sg13g2_nand3_1
XFILLER_56_966 VPWR VGND sg13g2_fill_2
XFILLER_16_808 VPWR VGND sg13g2_fill_2
XFILLER_27_112 VPWR VGND sg13g2_decap_8
XFILLER_28_635 VPWR VGND sg13g2_decap_4
XFILLER_82_262 VPWR VGND sg13g2_fill_2
XFILLER_27_167 VPWR VGND sg13g2_decap_4
X_09577_ _03693_ VPWR _03694_ VGND net1806 _03638_ sg13g2_o21ai_1
XFILLER_70_435 VPWR VGND sg13g2_decap_8
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_36_690 VPWR VGND sg13g2_decap_8
XFILLER_35_35 VPWR VGND sg13g2_decap_8
X_08528_ VPWR _02752_ _02751_ VGND sg13g2_inv_1
X_08459_ _02692_ _02684_ _02691_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_502 VPWR VGND sg13g2_decap_8
XFILLER_23_384 VPWR VGND sg13g2_fill_2
X_11470_ fpdiv.reg_b_out\[11\] fp16_res_pipe.x2\[11\] net1940 _01040_ VPWR VGND sg13g2_mux2_1
XFILLER_51_56 VPWR VGND sg13g2_decap_8
X_10421_ VPWR _04470_ _04469_ VGND sg13g2_inv_1
XFILLER_125_949 VPWR VGND sg13g2_decap_8
X_13140_ piso.tx_bit_counter\[4\] net3 _06890_ _06891_ VPWR VGND sg13g2_nor3_1
X_10352_ _04399_ _04401_ _04402_ VPWR VGND sg13g2_nor2_1
XFILLER_124_437 VPWR VGND sg13g2_fill_1
X_13071_ _06837_ _06838_ _06821_ _06839_ VPWR VGND sg13g2_nand3_1
X_12022_ _05871_ _05843_ _05839_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_756 VPWR VGND sg13g2_decap_8
X_10283_ _04322_ _04156_ _04352_ VPWR VGND sg13g2_nor2_1
XFILLER_104_172 VPWR VGND sg13g2_fill_1
XFILLER_120_665 VPWR VGND sg13g2_decap_8
XFILLER_116_82 VPWR VGND sg13g2_decap_8
XFILLER_66_719 VPWR VGND sg13g2_decap_8
X_13973_ VPWR _00524_ net25 VGND sg13g2_inv_1
XFILLER_74_730 VPWR VGND sg13g2_decap_4
X_12924_ _06698_ _06694_ _06697_ _06520_ net1949 VPWR VGND sg13g2_a22oi_1
XFILLER_46_421 VPWR VGND sg13g2_decap_4
XFILLER_47_999 VPWR VGND sg13g2_fill_2
XFILLER_47_988 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_18_156 VPWR VGND sg13g2_decap_8
X_12855_ _06634_ VPWR _06635_ VGND net1960 _06632_ sg13g2_o21ai_1
XFILLER_18_189 VPWR VGND sg13g2_decap_4
XFILLER_92_96 VPWR VGND sg13g2_fill_2
X_12786_ VGND VPWR _06570_ piso.tx_bit_counter\[3\] _06571_ piso.tx_bit_counter\[4\]
+ sg13g2_a21oi_1
X_11806_ _05621_ VPWR _05707_ VGND _05634_ _05641_ sg13g2_o21ai_1
X_14525_ _00326_ VGND VPWR _01061_ fpdiv.div_out\[0\] clknet_leaf_73_clk sg13g2_dfrbpq_1
XFILLER_42_671 VPWR VGND sg13g2_fill_2
XFILLER_42_660 VPWR VGND sg13g2_decap_8
XFILLER_15_896 VPWR VGND sg13g2_decap_8
XFILLER_30_822 VPWR VGND sg13g2_fill_1
X_11737_ _05638_ _05640_ _05641_ VPWR VGND sg13g2_nor2_1
XFILLER_41_181 VPWR VGND sg13g2_decap_4
XFILLER_30_833 VPWR VGND sg13g2_fill_2
XFILLER_30_855 VPWR VGND sg13g2_decap_8
XFILLER_30_866 VPWR VGND sg13g2_fill_1
X_14456_ _00257_ VGND VPWR _00995_ fpmul.seg_reg0.q\[41\] clknet_leaf_107_clk sg13g2_dfrbpq_1
X_11668_ fp16_sum_pipe.reg3en.q\[0\] _05573_ VPWR VGND sg13g2_inv_4
XFILLER_30_899 VPWR VGND sg13g2_decap_8
XFILLER_127_231 VPWR VGND sg13g2_decap_8
XFILLER_116_905 VPWR VGND sg13g2_decap_8
X_14387_ _00188_ VGND VPWR _00926_ div_result\[0\] clknet_leaf_75_clk sg13g2_dfrbpq_1
X_13407_ _07082_ net1721 instr\[13\] VPWR VGND sg13g2_nand2_1
X_10619_ _04619_ _04631_ _04632_ VPWR VGND sg13g2_nor2_1
X_11599_ _05421_ _05400_ _05418_ _05504_ VPWR VGND _05502_ sg13g2_nand4_1
Xplace1706 _02654_ net1706 VPWR VGND sg13g2_buf_2
Xplace1717 _06574_ net1717 VPWR VGND sg13g2_buf_2
X_13338_ _07041_ VPWR _00828_ VGND _07040_ net1726 sg13g2_o21ai_1
Xplace1728 _02574_ net1728 VPWR VGND sg13g2_buf_2
Xplace1739 _02726_ net1739 VPWR VGND sg13g2_buf_2
X_13269_ VGND VPWR net1676 _06987_ _00844_ _06988_ sg13g2_a21oi_1
XFILLER_111_621 VPWR VGND sg13g2_decap_8
XFILLER_69_513 VPWR VGND sg13g2_decap_8
XFILLER_110_120 VPWR VGND sg13g2_decap_4
X_07830_ _02126_ _02006_ acc_sub.exp_mant_logic0.b\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_97_866 VPWR VGND sg13g2_decap_8
XFILLER_99_1007 VPWR VGND sg13g2_decap_8
XFILLER_84_527 VPWR VGND sg13g2_fill_2
XFILLER_38_911 VPWR VGND sg13g2_decap_8
XFILLER_38_966 VPWR VGND sg13g2_decap_8
XFILLER_38_955 VPWR VGND sg13g2_fill_1
XFILLER_38_944 VPWR VGND sg13g2_decap_8
X_09500_ _03618_ acc_sub.x2\[0\] net1916 VPWR VGND sg13g2_nand2_1
X_07692_ _02000_ _01989_ net1792 VPWR VGND sg13g2_nand2_1
XFILLER_92_560 VPWR VGND sg13g2_decap_4
XFILLER_25_616 VPWR VGND sg13g2_decap_8
XFILLER_92_571 VPWR VGND sg13g2_decap_8
XFILLER_65_796 VPWR VGND sg13g2_decap_8
XFILLER_64_273 VPWR VGND sg13g2_fill_2
X_09431_ _03573_ _03450_ fp16_res_pipe.reg2en.q\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_52_468 VPWR VGND sg13g2_decap_4
X_09362_ VPWR _03512_ fp16_res_pipe.add_renorm0.mantisa\[8\] VGND sg13g2_inv_1
XFILLER_61_991 VPWR VGND sg13g2_fill_1
XFILLER_40_619 VPWR VGND sg13g2_fill_2
XFILLER_36_1013 VPWR VGND sg13g2_fill_1
XFILLER_33_682 VPWR VGND sg13g2_decap_8
X_08313_ _01362_ _02557_ _02558_ VPWR VGND sg13g2_nand2_1
XFILLER_21_800 VPWR VGND sg13g2_fill_1
XFILLER_21_811 VPWR VGND sg13g2_decap_8
X_09293_ VPWR _03447_ _03446_ VGND sg13g2_inv_1
XFILLER_21_855 VPWR VGND sg13g2_fill_1
X_08244_ _02496_ fp16_sum_pipe.exp_mant_logic0.b\[3\] _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[6\]
+ net1777 VPWR VGND sg13g2_a22oi_1
XFILLER_20_343 VPWR VGND sg13g2_decap_8
XFILLER_119_765 VPWR VGND sg13g2_decap_8
XFILLER_118_231 VPWR VGND sg13g2_decap_8
X_08175_ _01375_ _02432_ _02433_ VPWR VGND sg13g2_nand2_1
X_07126_ VPWR _01498_ acc_sub.seg_reg1.q\[20\] VGND sg13g2_inv_1
XFILLER_102_621 VPWR VGND sg13g2_decap_4
XFILLER_0_737 VPWR VGND sg13g2_fill_1
XFILLER_101_120 VPWR VGND sg13g2_decap_4
XFILLER_87_354 VPWR VGND sg13g2_fill_2
XFILLER_87_343 VPWR VGND sg13g2_fill_2
XFILLER_102_698 VPWR VGND sg13g2_fill_1
XFILLER_29_955 VPWR VGND sg13g2_decap_8
X_07959_ _02232_ VPWR _02233_ VGND _02206_ _02231_ sg13g2_o21ai_1
XFILLER_55_251 VPWR VGND sg13g2_fill_1
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_44_925 VPWR VGND sg13g2_fill_1
XFILLER_44_914 VPWR VGND sg13g2_decap_8
X_10970_ _04970_ net1710 _04681_ VPWR VGND sg13g2_nand2_1
X_09629_ net1804 VPWR _03746_ VGND _03675_ _03628_ sg13g2_o21ai_1
X_12640_ _06455_ VPWR _06456_ VGND net1851 _05339_ sg13g2_o21ai_1
XFILLER_62_33 VPWR VGND sg13g2_decap_8
XFILLER_24_671 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_50_clk clknet_5_22__leaf_clk clknet_leaf_50_clk VPWR VGND sg13g2_buf_8
X_12571_ _06387_ _06386_ _06383_ VPWR VGND sg13g2_nand2b_1
X_14310_ _00111_ VGND VPWR _00854_ sipo.bit_counter\[4\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_51_490 VPWR VGND sg13g2_decap_8
XFILLER_12_855 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
X_11522_ _05402_ _05425_ _05426_ _05427_ VPWR VGND sg13g2_nor3_2
XFILLER_127_0 VPWR VGND sg13g2_decap_8
X_11453_ VPWR _05378_ fpdiv.divider0.dividend\[7\] VGND sg13g2_inv_1
X_14241_ _00042_ VGND VPWR _00792_ instr\[6\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_14172_ VPWR _00723_ net105 VGND sg13g2_inv_1
X_10404_ VPWR _04454_ _04453_ VGND sg13g2_inv_1
XFILLER_125_746 VPWR VGND sg13g2_decap_8
X_13123_ VGND VPWR _06877_ _06792_ _06868_ sg13g2_or2_1
X_11384_ _05332_ _05333_ _05331_ _05334_ VPWR VGND sg13g2_nand3_1
XFILLER_127_70 VPWR VGND sg13g2_decap_8
XFILLER_124_245 VPWR VGND sg13g2_decap_8
XFILLER_106_971 VPWR VGND sg13g2_decap_8
XFILLER_3_553 VPWR VGND sg13g2_decap_8
XFILLER_11_70 VPWR VGND sg13g2_decap_8
X_10335_ _04386_ _04384_ VPWR VGND sg13g2_inv_2
X_13054_ fpmul.seg_reg0.q\[49\] fpmul.seg_reg0.q\[48\] fpmul.seg_reg0.q\[47\] fpmul.seg_reg0.q\[46\]
+ _06822_ VPWR VGND sg13g2_nor4_1
X_10266_ _04336_ _04224_ net1745 VPWR VGND sg13g2_nand2_1
XFILLER_121_952 VPWR VGND sg13g2_decap_8
XFILLER_94_803 VPWR VGND sg13g2_decap_8
XFILLER_78_343 VPWR VGND sg13g2_decap_8
X_12005_ _05859_ _05825_ _05858_ VPWR VGND sg13g2_xnor2_1
XFILLER_120_451 VPWR VGND sg13g2_fill_1
XFILLER_94_836 VPWR VGND sg13g2_decap_8
XFILLER_79_888 VPWR VGND sg13g2_decap_8
XFILLER_78_387 VPWR VGND sg13g2_fill_2
XFILLER_78_365 VPWR VGND sg13g2_decap_4
XFILLER_4_1000 VPWR VGND sg13g2_decap_8
X_10197_ _04274_ net1636 _04271_ VPWR VGND sg13g2_nand2b_1
XFILLER_66_538 VPWR VGND sg13g2_decap_4
XFILLER_16_7 VPWR VGND sg13g2_decap_8
X_13956_ VPWR _00507_ net92 VGND sg13g2_inv_1
XFILLER_81_508 VPWR VGND sg13g2_fill_2
XFILLER_74_560 VPWR VGND sg13g2_fill_1
XFILLER_62_700 VPWR VGND sg13g2_decap_4
X_12907_ _00011_ net1731 net1702 _06682_ VPWR VGND sg13g2_nand3_1
XFILLER_62_722 VPWR VGND sg13g2_fill_2
XFILLER_35_925 VPWR VGND sg13g2_decap_8
X_13887_ VPWR _00438_ net49 VGND sg13g2_inv_1
X_12838_ _06618_ _06617_ net1922 _06619_ VPWR VGND sg13g2_a21o_2
XFILLER_15_660 VPWR VGND sg13g2_decap_8
X_12769_ _00008_ _00007_ _00006_ _00005_ _06554_ VPWR VGND sg13g2_nor4_1
XFILLER_14_181 VPWR VGND sg13g2_fill_1
X_14508_ _00309_ VGND VPWR _01044_ fpdiv.reg_b_out\[15\] clknet_leaf_91_clk sg13g2_dfrbpq_1
X_14439_ _00240_ VGND VPWR _00978_ fpmul.seg_reg0.q\[24\] clknet_leaf_105_clk sg13g2_dfrbpq_1
XFILLER_7_881 VPWR VGND sg13g2_decap_8
XFILLER_116_779 VPWR VGND sg13g2_decap_8
XFILLER_115_245 VPWR VGND sg13g2_decap_8
XFILLER_104_908 VPWR VGND sg13g2_decap_8
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_09980_ fp16_res_pipe.exp_mant_logic0.a\[10\] fp16_res_pipe.exp_mant_logic0.a\[9\]
+ fp16_res_pipe.exp_mant_logic0.a\[8\] fp16_res_pipe.exp_mant_logic0.a\[7\] _04069_
+ VPWR VGND sg13g2_nor4_1
X_08931_ _03116_ _03117_ _03115_ _03118_ VPWR VGND sg13g2_nand3_1
XFILLER_103_429 VPWR VGND sg13g2_decap_8
XFILLER_69_310 VPWR VGND sg13g2_decap_8
X_08862_ _03049_ _03010_ _02971_ VPWR VGND sg13g2_nand2_1
XFILLER_97_652 VPWR VGND sg13g2_fill_1
XFILLER_112_985 VPWR VGND sg13g2_decap_8
X_07813_ _01414_ _02109_ _02110_ VPWR VGND sg13g2_nand2_1
XFILLER_84_302 VPWR VGND sg13g2_decap_8
XFILLER_29_207 VPWR VGND sg13g2_decap_8
XFILLER_29_218 VPWR VGND sg13g2_fill_2
XFILLER_123_28 VPWR VGND sg13g2_decap_8
X_07744_ _01753_ _02048_ _02049_ VPWR VGND sg13g2_nor2_1
XFILLER_38_763 VPWR VGND sg13g2_fill_1
X_07675_ _01985_ _01984_ net1641 VPWR VGND sg13g2_nand2_1
XFILLER_93_891 VPWR VGND sg13g2_decap_8
XFILLER_53_722 VPWR VGND sg13g2_decap_8
XFILLER_25_424 VPWR VGND sg13g2_decap_8
XFILLER_26_947 VPWR VGND sg13g2_decap_8
XFILLER_53_766 VPWR VGND sg13g2_fill_2
X_09414_ _03558_ net1675 _03489_ VPWR VGND sg13g2_nand2_1
XFILLER_80_574 VPWR VGND sg13g2_decap_8
XFILLER_41_928 VPWR VGND sg13g2_decap_8
XFILLER_40_416 VPWR VGND sg13g2_decap_8
XFILLER_12_118 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_32_clk clknet_5_17__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
X_09345_ _03497_ _03438_ _03496_ _03486_ _03374_ VPWR VGND sg13g2_a22oi_1
X_09276_ _03429_ VPWR _03430_ VGND _03397_ _03427_ sg13g2_o21ai_1
XFILLER_32_14 VPWR VGND sg13g2_decap_8
XFILLER_120_7 VPWR VGND sg13g2_decap_8
X_08227_ _02481_ net1691 net1842 VPWR VGND sg13g2_nand2_1
XFILLER_119_551 VPWR VGND sg13g2_decap_8
XFILLER_5_829 VPWR VGND sg13g2_decap_8
XFILLER_119_595 VPWR VGND sg13g2_decap_8
XFILLER_119_584 VPWR VGND sg13g2_decap_4
XFILLER_107_724 VPWR VGND sg13g2_decap_8
XFILLER_4_317 VPWR VGND sg13g2_fill_2
X_08158_ _02418_ _02417_ net1639 VPWR VGND sg13g2_nand2_1
X_08089_ _02355_ fp16_sum_pipe.exp_mant_logic0.a\[6\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[9\]
+ net1776 VPWR VGND sg13g2_a22oi_1
XFILLER_122_749 VPWR VGND sg13g2_decap_8
XFILLER_79_118 VPWR VGND sg13g2_decap_8
XFILLER_0_512 VPWR VGND sg13g2_decap_8
X_10120_ _03609_ _04140_ _04203_ VPWR VGND sg13g2_nor2_1
XFILLER_121_259 VPWR VGND sg13g2_decap_8
XFILLER_88_630 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_99_clk clknet_5_15__leaf_clk clknet_leaf_99_clk VPWR VGND sg13g2_buf_8
XFILLER_0_556 VPWR VGND sg13g2_decap_8
X_10051_ VPWR _04139_ _04138_ VGND sg13g2_inv_1
XFILLER_103_974 VPWR VGND sg13g2_decap_8
XFILLER_57_11 VPWR VGND sg13g2_fill_2
X_13810_ VPWR _00361_ net77 VGND sg13g2_inv_1
X_14790_ _00591_ VGND VPWR _01314_ acc_sum.exp_mant_logic0.a\[3\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
XFILLER_91_839 VPWR VGND sg13g2_decap_8
X_13741_ VPWR _00292_ net86 VGND sg13g2_inv_1
XFILLER_16_424 VPWR VGND sg13g2_fill_2
XFILLER_17_947 VPWR VGND sg13g2_decap_8
X_10953_ fp16_res_pipe.seg_reg1.q\[21\] _04957_ _04958_ _04959_ VPWR VGND sg13g2_nor3_1
XFILLER_83_390 VPWR VGND sg13g2_fill_2
XFILLER_73_43 VPWR VGND sg13g2_fill_1
XFILLER_44_744 VPWR VGND sg13g2_fill_2
XFILLER_43_221 VPWR VGND sg13g2_decap_8
X_13672_ VPWR _00223_ net122 VGND sg13g2_inv_1
XFILLER_73_87 VPWR VGND sg13g2_fill_2
X_10884_ _04737_ _04894_ _04893_ _04895_ VPWR VGND sg13g2_nand3_1
XFILLER_25_980 VPWR VGND sg13g2_decap_8
X_12623_ _06439_ _05342_ net1852 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_23_clk clknet_5_19__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_31_427 VPWR VGND sg13g2_decap_8
X_12554_ _06370_ VPWR _00941_ VGND _06354_ _06369_ sg13g2_o21ai_1
XFILLER_8_656 VPWR VGND sg13g2_decap_8
XFILLER_8_634 VPWR VGND sg13g2_decap_8
X_11505_ _05410_ net1840 fp16_sum_pipe.add_renorm0.mantisa\[3\] VPWR VGND sg13g2_nand2_1
X_12485_ _06323_ _06321_ _06322_ VPWR VGND sg13g2_xnor2_1
X_14224_ _00025_ VGND VPWR _00775_ sipo.shift_reg\[5\] clknet_leaf_14_clk sg13g2_dfrbpq_1
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_11_184 VPWR VGND sg13g2_decap_8
X_11436_ _05367_ acc_sub.x2\[9\] VPWR VGND sg13g2_inv_2
X_14155_ VPWR _00706_ net130 VGND sg13g2_inv_1
X_11367_ _01075_ _05317_ _05318_ VPWR VGND sg13g2_nand2_1
X_14086_ VPWR _00637_ net89 VGND sg13g2_inv_1
X_13106_ VGND VPWR _06774_ _06856_ _06864_ _06835_ sg13g2_a21oi_1
XFILLER_4_895 VPWR VGND sg13g2_decap_8
X_10318_ _04376_ VPWR _01182_ VGND net1919 _04012_ sg13g2_o21ai_1
X_13037_ VPWR _06805_ _06804_ VGND sg13g2_inv_1
XFILLER_67_803 VPWR VGND sg13g2_fill_1
XFILLER_39_505 VPWR VGND sg13g2_fill_2
X_10249_ _04320_ _04158_ fp16_res_pipe.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_78_184 VPWR VGND sg13g2_decap_8
XFILLER_66_335 VPWR VGND sg13g2_decap_8
XFILLER_39_549 VPWR VGND sg13g2_decap_8
XFILLER_120_292 VPWR VGND sg13g2_decap_4
XFILLER_82_817 VPWR VGND sg13g2_decap_4
XFILLER_81_327 VPWR VGND sg13g2_decap_8
XFILLER_19_262 VPWR VGND sg13g2_decap_8
X_13939_ VPWR _00490_ net26 VGND sg13g2_inv_1
XFILLER_34_243 VPWR VGND sg13g2_fill_1
X_07460_ acc_sub.exp_mant_logic0.b\[13\] _01727_ _01783_ VPWR VGND sg13g2_nor2_1
XFILLER_16_980 VPWR VGND sg13g2_decap_8
X_07391_ _01736_ net1894 acc\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_72_1010 VPWR VGND sg13g2_decap_4
XFILLER_50_736 VPWR VGND sg13g2_decap_8
X_09130_ net1785 _03308_ _03309_ _03310_ VPWR VGND sg13g2_nor3_1
Xclkbuf_leaf_14_clk clknet_5_4__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_09061_ _03198_ _03245_ _03246_ VPWR VGND sg13g2_nor2_1
X_08012_ _02277_ VPWR _02278_ VGND _02219_ _02214_ sg13g2_o21ai_1
XFILLER_118_28 VPWR VGND sg13g2_decap_8
XFILLER_116_521 VPWR VGND sg13g2_decap_8
XFILLER_89_438 VPWR VGND sg13g2_decap_4
XFILLER_1_309 VPWR VGND sg13g2_decap_4
X_08914_ _03097_ _03100_ _03101_ VPWR VGND sg13g2_nor2_1
X_09894_ fp16_res_pipe.exp_mant_logic0.b\[14\] net1765 _03991_ VPWR VGND sg13g2_nor2_1
X_08845_ _03023_ _03027_ _03031_ _03032_ VPWR VGND sg13g2_nor3_1
XFILLER_112_782 VPWR VGND sg13g2_decap_8
XFILLER_100_944 VPWR VGND sg13g2_decap_8
XFILLER_58_847 VPWR VGND sg13g2_fill_2
X_08776_ _02964_ acc\[0\] net1896 VPWR VGND sg13g2_nand2_1
XFILLER_57_368 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
X_07727_ _01747_ _01977_ _02033_ VPWR VGND sg13g2_nor2_1
XFILLER_72_338 VPWR VGND sg13g2_fill_2
XFILLER_72_305 VPWR VGND sg13g2_fill_1
XFILLER_25_210 VPWR VGND sg13g2_fill_1
X_07658_ _01969_ acc_sub.exp_mant_logic0.a\[4\] net1651 net1685 acc_sub.exp_mant_logic0.a\[3\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_13_405 VPWR VGND sg13g2_fill_1
XFILLER_25_276 VPWR VGND sg13g2_fill_1
XFILLER_26_799 VPWR VGND sg13g2_decap_8
X_07589_ _01903_ _01873_ _01902_ VPWR VGND sg13g2_xnor2_1
XFILLER_80_382 VPWR VGND sg13g2_decap_8
Xclkbuf_4_8_0_clk clknet_0_clk clknet_4_8_0_clk VPWR VGND sg13g2_buf_8
XFILLER_53_596 VPWR VGND sg13g2_fill_2
XFILLER_43_35 VPWR VGND sg13g2_decap_8
XFILLER_41_747 VPWR VGND sg13g2_decap_4
X_09328_ _03481_ _03480_ _03365_ VPWR VGND sg13g2_nand2_1
XFILLER_22_961 VPWR VGND sg13g2_decap_8
X_09259_ _03413_ _03412_ fp16_res_pipe.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_126_329 VPWR VGND sg13g2_decap_8
XFILLER_119_370 VPWR VGND sg13g2_decap_8
X_12270_ VGND VPWR _06101_ _06094_ _06116_ _06115_ sg13g2_a21oi_1
XFILLER_104_2 VPWR VGND sg13g2_fill_1
X_11221_ _05187_ _05178_ _05186_ VPWR VGND sg13g2_nand2_1
XFILLER_4_147 VPWR VGND sg13g2_decap_8
X_11152_ _05122_ _05121_ VPWR VGND sg13g2_inv_2
XFILLER_1_843 VPWR VGND sg13g2_decap_8
X_10103_ VGND VPWR _04165_ net1828 _04187_ _04186_ sg13g2_a21oi_1
XFILLER_110_708 VPWR VGND sg13g2_fill_2
XFILLER_89_972 VPWR VGND sg13g2_decap_8
XFILLER_76_600 VPWR VGND sg13g2_decap_8
X_11083_ _05059_ _04993_ acc_sum.seg_reg0.q\[26\] VPWR VGND sg13g2_nand2_1
X_14911_ _00712_ VGND VPWR _01431_ acc_sub.op_sign_logic0.mantisa_a\[10\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_1
XFILLER_49_858 VPWR VGND sg13g2_fill_1
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_0_386 VPWR VGND sg13g2_decap_8
X_10034_ VPWR _04122_ _04121_ VGND sg13g2_inv_1
XFILLER_48_346 VPWR VGND sg13g2_fill_1
X_14842_ _00643_ VGND VPWR _01366_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[4\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
XFILLER_57_891 VPWR VGND sg13g2_fill_1
X_14773_ _00574_ VGND VPWR _01297_ acc_sub.y\[2\] clknet_leaf_46_clk sg13g2_dfrbpq_1
XFILLER_63_349 VPWR VGND sg13g2_decap_8
X_11985_ _05839_ _05837_ _05838_ VPWR VGND sg13g2_xnor2_1
X_13724_ VPWR _00275_ net137 VGND sg13g2_inv_1
XFILLER_72_861 VPWR VGND sg13g2_fill_1
XFILLER_44_574 VPWR VGND sg13g2_decap_8
XFILLER_44_552 VPWR VGND sg13g2_decap_4
XFILLER_16_243 VPWR VGND sg13g2_decap_4
X_10936_ _04740_ _04809_ _04943_ VPWR VGND sg13g2_nor2_1
XFILLER_32_714 VPWR VGND sg13g2_fill_2
X_13655_ VPWR _00206_ net68 VGND sg13g2_inv_1
X_10867_ _04860_ _04878_ _04879_ VPWR VGND sg13g2_nor2_1
XFILLER_31_224 VPWR VGND sg13g2_decap_8
X_12606_ _06422_ _06421_ _05348_ VPWR VGND sg13g2_nand2_1
XFILLER_13_961 VPWR VGND sg13g2_decap_8
XFILLER_83_7 VPWR VGND sg13g2_decap_4
X_13586_ VPWR _00137_ net121 VGND sg13g2_inv_1
X_10798_ _04810_ _04809_ _04740_ VPWR VGND sg13g2_nand2_1
XFILLER_31_279 VPWR VGND sg13g2_fill_2
X_12537_ _02648_ _06354_ VPWR VGND sg13g2_inv_4
XFILLER_9_976 VPWR VGND sg13g2_decap_8
XFILLER_117_329 VPWR VGND sg13g2_fill_2
XFILLER_117_318 VPWR VGND sg13g2_decap_8
X_12468_ _06310_ _06309_ _06056_ VPWR VGND sg13g2_nand2_1
XFILLER_8_497 VPWR VGND sg13g2_decap_8
XFILLER_126_841 VPWR VGND sg13g2_decap_8
X_14207_ VPWR _00758_ net106 VGND sg13g2_inv_1
X_11419_ fpdiv.reg_a_out\[15\] net1942 _05356_ VPWR VGND sg13g2_nor2_1
XFILLER_125_373 VPWR VGND sg13g2_decap_4
XFILLER_113_524 VPWR VGND sg13g2_fill_1
XFILLER_113_513 VPWR VGND sg13g2_fill_2
X_14138_ VPWR _00689_ net114 VGND sg13g2_inv_1
X_12399_ _06245_ _06244_ _06209_ VPWR VGND sg13g2_nand2_1
XFILLER_87_909 VPWR VGND sg13g2_decap_8
X_14069_ VPWR _00620_ net95 VGND sg13g2_inv_1
XFILLER_98_257 VPWR VGND sg13g2_decap_8
XFILLER_67_600 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_3_clk clknet_5_5__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
XFILLER_100_229 VPWR VGND sg13g2_fill_1
XFILLER_95_953 VPWR VGND sg13g2_decap_8
XFILLER_39_313 VPWR VGND sg13g2_decap_8
X_08630_ VGND VPWR _02851_ _02778_ _02852_ _02777_ sg13g2_a21oi_1
XFILLER_82_636 VPWR VGND sg13g2_fill_2
XFILLER_82_625 VPWR VGND sg13g2_decap_8
X_08561_ VGND VPWR _02769_ _02782_ _02785_ _02784_ sg13g2_a21oi_1
XFILLER_66_198 VPWR VGND sg13g2_decap_4
X_08492_ _02719_ _02692_ fpdiv.divider0.divisor_reg\[4\] VPWR VGND sg13g2_nand2_1
X_07512_ VPWR _01834_ _01796_ VGND sg13g2_inv_1
XFILLER_81_179 VPWR VGND sg13g2_decap_8
X_07443_ VPWR _01772_ fpdiv.divider0.divisor_reg\[5\] VGND sg13g2_inv_1
Xfanout17 net18 net17 VPWR VGND sg13g2_buf_2
Xfanout28 net31 net28 VPWR VGND sg13g2_buf_2
XFILLER_22_213 VPWR VGND sg13g2_fill_1
Xfanout39 net72 net39 VPWR VGND sg13g2_buf_2
XFILLER_50_555 VPWR VGND sg13g2_decap_8
XFILLER_22_246 VPWR VGND sg13g2_decap_8
XFILLER_23_769 VPWR VGND sg13g2_decap_8
X_09113_ _03294_ acc_sub.y\[9\] VPWR VGND sg13g2_inv_2
X_07374_ VGND VPWR _01723_ net1893 _01467_ _01724_ sg13g2_a21oi_1
XFILLER_13_49 VPWR VGND sg13g2_decap_8
XFILLER_31_791 VPWR VGND sg13g2_decap_8
XFILLER_117_830 VPWR VGND sg13g2_decap_8
X_09044_ VPWR _03230_ _03229_ VGND sg13g2_inv_1
XFILLER_116_373 VPWR VGND sg13g2_fill_2
XFILLER_89_279 VPWR VGND sg13g2_fill_2
XFILLER_89_268 VPWR VGND sg13g2_decap_8
X_09946_ VPWR _04042_ _03994_ VGND sg13g2_inv_1
XFILLER_86_931 VPWR VGND sg13g2_decap_8
XFILLER_38_35 VPWR VGND sg13g2_decap_8
X_09877_ acc_sum.y\[2\] _03765_ net1820 _01227_ VPWR VGND sg13g2_mux2_1
XFILLER_97_290 VPWR VGND sg13g2_fill_2
X_08759_ _02952_ VPWR _01317_ VGND net1899 _02951_ sg13g2_o21ai_1
XFILLER_72_124 VPWR VGND sg13g2_decap_8
XFILLER_54_872 VPWR VGND sg13g2_decap_8
XFILLER_54_56 VPWR VGND sg13g2_fill_1
X_11770_ _05674_ _05652_ _05673_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_574 VPWR VGND sg13g2_decap_8
XFILLER_54_89 VPWR VGND sg13g2_decap_8
XFILLER_41_533 VPWR VGND sg13g2_decap_8
X_10721_ _04681_ _04672_ _04642_ _04675_ _04734_ VPWR VGND sg13g2_nor4_1
X_13440_ _07099_ net1751 sipo.shift_reg\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_41_566 VPWR VGND sg13g2_decap_4
XFILLER_9_206 VPWR VGND sg13g2_fill_2
XFILLER_14_758 VPWR VGND sg13g2_fill_1
XFILLER_110_95 VPWR VGND sg13g2_decap_8
XFILLER_110_84 VPWR VGND sg13g2_decap_4
X_10652_ _04665_ _04660_ _04664_ VPWR VGND sg13g2_nand2_2
X_13371_ _07061_ VPWR _00815_ VGND _05359_ net1694 sg13g2_o21ai_1
X_10583_ _04604_ VPWR _01145_ VGND net1932 _02264_ sg13g2_o21ai_1
XFILLER_126_126 VPWR VGND sg13g2_decap_8
XFILLER_70_88 VPWR VGND sg13g2_fill_1
X_12322_ _06167_ _06160_ _06168_ VPWR VGND sg13g2_xor2_1
XFILLER_6_913 VPWR VGND sg13g2_decap_8
XFILLER_10_975 VPWR VGND sg13g2_decap_8
X_12253_ _06075_ _06071_ _06099_ VPWR VGND sg13g2_nor2b_1
XFILLER_107_351 VPWR VGND sg13g2_decap_4
X_11204_ _05171_ net1635 _05170_ VPWR VGND sg13g2_nand2_1
XFILLER_5_478 VPWR VGND sg13g2_decap_8
XFILLER_123_855 VPWR VGND sg13g2_decap_8
XFILLER_122_310 VPWR VGND sg13g2_fill_1
XFILLER_79_97 VPWR VGND sg13g2_decap_8
X_12184_ VPWR _06030_ _06029_ VGND sg13g2_inv_1
XFILLER_122_354 VPWR VGND sg13g2_fill_1
X_11135_ _05098_ _05101_ _05104_ _05105_ VPWR VGND sg13g2_nor3_1
XFILLER_49_600 VPWR VGND sg13g2_decap_8
XFILLER_122_387 VPWR VGND sg13g2_decap_4
XFILLER_110_538 VPWR VGND sg13g2_fill_2
X_11066_ VGND VPWR _05042_ _02937_ _05044_ _04993_ sg13g2_a21oi_1
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_95_63 VPWR VGND sg13g2_fill_2
XFILLER_76_452 VPWR VGND sg13g2_fill_1
XFILLER_76_441 VPWR VGND sg13g2_fill_1
X_10017_ _04090_ _04104_ _04105_ VPWR VGND sg13g2_nor2_2
XFILLER_63_102 VPWR VGND sg13g2_fill_2
XFILLER_36_316 VPWR VGND sg13g2_decap_4
X_14825_ _00626_ VGND VPWR _01349_ fpdiv.divider0.remainder_reg\[4\] clknet_leaf_70_clk
+ sg13g2_dfrbpq_2
XFILLER_92_967 VPWR VGND sg13g2_decap_8
XFILLER_64_669 VPWR VGND sg13g2_decap_4
XFILLER_63_124 VPWR VGND sg13g2_fill_1
X_14756_ _00557_ VGND VPWR _01280_ acc_sum.exp_mant_logic0.b\[1\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_91_499 VPWR VGND sg13g2_decap_4
X_13707_ VPWR _00258_ net64 VGND sg13g2_inv_1
X_11968_ _05822_ VPWR _00978_ VGND net1884 _05821_ sg13g2_o21ai_1
XFILLER_17_585 VPWR VGND sg13g2_fill_1
XFILLER_32_533 VPWR VGND sg13g2_fill_1
X_11899_ _05780_ net1877 fpmul.reg_a_out\[11\] VPWR VGND sg13g2_nand2_1
X_10919_ _04928_ _04772_ fp16_res_pipe.y\[11\] VPWR VGND sg13g2_nand2_1
X_14687_ _00488_ VGND VPWR _01215_ fp16_res_pipe.seg_reg0.q\[24\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_1
XFILLER_32_544 VPWR VGND sg13g2_decap_8
XFILLER_81_4 VPWR VGND sg13g2_fill_2
X_13638_ VPWR _00189_ net124 VGND sg13g2_inv_1
X_13569_ VPWR _00120_ net34 VGND sg13g2_inv_1
XFILLER_118_638 VPWR VGND sg13g2_fill_2
XFILLER_117_126 VPWR VGND sg13g2_decap_8
XFILLER_9_795 VPWR VGND sg13g2_decap_8
XFILLER_114_811 VPWR VGND sg13g2_decap_8
XFILLER_119_1010 VPWR VGND sg13g2_decap_4
XFILLER_99_555 VPWR VGND sg13g2_fill_2
XFILLER_5_990 VPWR VGND sg13g2_decap_8
XFILLER_114_888 VPWR VGND sg13g2_decap_8
X_09800_ _03648_ VPWR _03914_ VGND _03873_ _03913_ sg13g2_o21ai_1
XFILLER_101_505 VPWR VGND sg13g2_fill_2
XFILLER_99_566 VPWR VGND sg13g2_fill_2
X_07992_ VPWR _02259_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[10\] VGND sg13g2_inv_1
X_09731_ _03845_ _03846_ _03847_ VPWR VGND sg13g2_nor2_1
XFILLER_68_920 VPWR VGND sg13g2_fill_1
XFILLER_67_441 VPWR VGND sg13g2_decap_4
X_09662_ VGND VPWR _03778_ _03779_ _03776_ _03740_ sg13g2_a21oi_2
XFILLER_68_997 VPWR VGND sg13g2_fill_1
XFILLER_68_986 VPWR VGND sg13g2_decap_8
XFILLER_67_485 VPWR VGND sg13g2_decap_8
XFILLER_67_463 VPWR VGND sg13g2_decap_8
XFILLER_55_614 VPWR VGND sg13g2_fill_1
XFILLER_39_154 VPWR VGND sg13g2_decap_4
X_09593_ _03710_ _03709_ VPWR VGND sg13g2_inv_2
X_08613_ _02836_ _02835_ _02812_ VPWR VGND sg13g2_nand2b_1
XFILLER_83_967 VPWR VGND sg13g2_decap_8
X_08544_ VPWR VGND _02767_ _02752_ _02759_ _02748_ _02768_ _02753_ sg13g2_a221oi_1
XFILLER_82_455 VPWR VGND sg13g2_fill_1
X_08475_ _02705_ VPWR _01354_ VGND net1705 _02704_ sg13g2_o21ai_1
X_07426_ VPWR _01760_ fpdiv.divider0.divisor_reg\[10\] VGND sg13g2_inv_1
XFILLER_51_886 VPWR VGND sg13g2_decap_8
XFILLER_50_374 VPWR VGND sg13g2_fill_1
X_07357_ _01714_ net1799 acc_sub.seg_reg0.q\[27\] VPWR VGND sg13g2_nand2_1
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_14 VPWR VGND sg13g2_decap_8
X_07288_ _01655_ VPWR _01484_ VGND acc_sub.reg2en.q\[0\] _01647_ sg13g2_o21ai_1
X_09027_ VGND VPWR _03193_ _03211_ _03213_ _03212_ sg13g2_a21oi_1
XFILLER_3_938 VPWR VGND sg13g2_decap_8
XFILLER_105_844 VPWR VGND sg13g2_decap_8
XFILLER_2_437 VPWR VGND sg13g2_decap_8
XFILLER_105_888 VPWR VGND sg13g2_decap_8
XFILLER_104_365 VPWR VGND sg13g2_decap_8
XFILLER_104_376 VPWR VGND sg13g2_fill_2
XFILLER_77_216 VPWR VGND sg13g2_decap_8
XFILLER_59_931 VPWR VGND sg13g2_fill_2
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_120_869 VPWR VGND sg13g2_decap_8
XFILLER_86_750 VPWR VGND sg13g2_fill_1
XFILLER_59_953 VPWR VGND sg13g2_decap_4
XFILLER_58_452 VPWR VGND sg13g2_fill_2
XFILLER_58_441 VPWR VGND sg13g2_decap_8
X_09929_ _04021_ _04025_ _04026_ VPWR VGND sg13g2_nor2_1
XFILLER_19_806 VPWR VGND sg13g2_fill_1
X_12940_ _06713_ _06712_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_59_997 VPWR VGND sg13g2_fill_2
XFILLER_59_986 VPWR VGND sg13g2_decap_8
XFILLER_18_316 VPWR VGND sg13g2_fill_1
XFILLER_19_839 VPWR VGND sg13g2_decap_8
XFILLER_74_967 VPWR VGND sg13g2_fill_2
X_12871_ _00014_ net1730 net1701 _06649_ VPWR VGND sg13g2_nand3_1
XFILLER_65_99 VPWR VGND sg13g2_fill_2
XFILLER_65_88 VPWR VGND sg13g2_fill_2
XFILLER_61_606 VPWR VGND sg13g2_fill_2
XFILLER_45_168 VPWR VGND sg13g2_decap_8
X_11822_ _05648_ VPWR _05722_ VGND _05642_ _05721_ sg13g2_o21ai_1
X_14610_ _00411_ VGND VPWR _01142_ fp16_sum_pipe.exp_mant_logic0.a\[5\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_2
XFILLER_92_1013 VPWR VGND sg13g2_fill_1
XFILLER_92_1002 VPWR VGND sg13g2_decap_8
XFILLER_60_127 VPWR VGND sg13g2_decap_4
XFILLER_42_831 VPWR VGND sg13g2_decap_8
XFILLER_26_360 VPWR VGND sg13g2_decap_8
XFILLER_27_883 VPWR VGND sg13g2_decap_8
XFILLER_81_54 VPWR VGND sg13g2_fill_1
XFILLER_81_43 VPWR VGND sg13g2_decap_8
XFILLER_81_32 VPWR VGND sg13g2_fill_1
X_14541_ _00342_ VGND VPWR _01077_ acc_sum.op_sign_logic0.mantisa_b\[4\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
XFILLER_26_393 VPWR VGND sg13g2_fill_1
X_11753_ _05657_ _04465_ fp16_sum_pipe.add_renorm0.exp\[3\] VPWR VGND sg13g2_nand2_1
X_14472_ _00273_ VGND VPWR _01011_ fpdiv.divider0.counter\[2\] clknet_leaf_73_clk
+ sg13g2_dfrbpq_1
X_10704_ _04637_ _04716_ _04717_ VPWR VGND sg13g2_nor2_1
X_13423_ _07090_ VPWR _00792_ VGND _06999_ net1719 sg13g2_o21ai_1
XFILLER_14_70 VPWR VGND sg13g2_decap_8
XFILLER_127_413 VPWR VGND sg13g2_fill_2
Xclkload109 clkload109/Y clknet_leaf_70_clk VPWR VGND sg13g2_inv_2
X_13354_ _07051_ net1723 fp16_res_pipe.x2\[3\] VPWR VGND sg13g2_nand2_1
X_12305_ _06151_ _06150_ _06134_ VPWR VGND sg13g2_xnor2_1
X_10566_ _04596_ fp16_sum_pipe.seg_reg0.q\[22\] net1845 VPWR VGND sg13g2_nand2_1
X_13285_ VPWR VGND acc_sub.y\[6\] _07000_ _02578_ net1728 _07001_ acc_sum.y\[6\] sg13g2_a221oi_1
XFILLER_5_264 VPWR VGND sg13g2_fill_1
X_10497_ _04541_ VPWR _04542_ VGND _04537_ _04540_ sg13g2_o21ai_1
XFILLER_108_682 VPWR VGND sg13g2_decap_8
X_12236_ _06063_ _06066_ _06082_ VPWR VGND sg13g2_nor2_1
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_6_798 VPWR VGND sg13g2_fill_2
XFILLER_5_297 VPWR VGND sg13g2_decap_8
XFILLER_30_91 VPWR VGND sg13g2_fill_2
XFILLER_123_663 VPWR VGND sg13g2_fill_1
XFILLER_123_652 VPWR VGND sg13g2_decap_4
XFILLER_122_140 VPWR VGND sg13g2_decap_8
XFILLER_111_803 VPWR VGND sg13g2_decap_8
X_12167_ _06013_ _06012_ _05980_ VPWR VGND sg13g2_nand2_1
XFILLER_123_685 VPWR VGND sg13g2_decap_4
XFILLER_110_302 VPWR VGND sg13g2_decap_8
XFILLER_96_547 VPWR VGND sg13g2_decap_8
X_11118_ _05009_ VPWR _05088_ VGND _05007_ _05087_ sg13g2_o21ai_1
XFILLER_2_982 VPWR VGND sg13g2_decap_8
XFILLER_96_558 VPWR VGND sg13g2_fill_2
X_12098_ VPWR _05944_ _05905_ VGND sg13g2_inv_1
XFILLER_49_430 VPWR VGND sg13g2_fill_2
XFILLER_1_492 VPWR VGND sg13g2_decap_8
XFILLER_77_794 VPWR VGND sg13g2_decap_8
X_11049_ _05028_ _05026_ acc_sum.exp_mant_logic0.a\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_92_753 VPWR VGND sg13g2_decap_4
XFILLER_49_496 VPWR VGND sg13g2_fill_1
X_14808_ _00609_ VGND VPWR _01332_ acc_sum.add_renorm0.exp\[5\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
XFILLER_52_628 VPWR VGND sg13g2_decap_8
XFILLER_33_820 VPWR VGND sg13g2_decap_4
XFILLER_17_360 VPWR VGND sg13g2_decap_8
XFILLER_17_371 VPWR VGND sg13g2_fill_1
XFILLER_33_853 VPWR VGND sg13g2_fill_1
X_14739_ _00540_ VGND VPWR _01267_ fp16_res_pipe.add_renorm0.mantisa\[2\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_2
XFILLER_32_330 VPWR VGND sg13g2_fill_1
XFILLER_33_897 VPWR VGND sg13g2_decap_8
X_08260_ _02471_ _02396_ _02510_ VPWR VGND sg13g2_nor2_1
XFILLER_32_374 VPWR VGND sg13g2_decap_8
X_07211_ _01500_ _01502_ _01583_ VPWR VGND sg13g2_nor2_1
X_08191_ _02445_ _02446_ _02447_ _02448_ VPWR VGND sg13g2_nor3_1
XFILLER_20_536 VPWR VGND sg13g2_fill_1
XFILLER_20_547 VPWR VGND sg13g2_fill_2
XFILLER_119_947 VPWR VGND sg13g2_decap_8
XFILLER_118_424 VPWR VGND sg13g2_decap_8
X_07142_ VPWR _01514_ _01513_ VGND sg13g2_inv_1
XFILLER_72_0 VPWR VGND sg13g2_fill_2
XFILLER_9_592 VPWR VGND sg13g2_decap_8
XFILLER_10_28 VPWR VGND sg13g2_decap_8
XFILLER_126_28 VPWR VGND sg13g2_decap_8
XFILLER_113_140 VPWR VGND sg13g2_decap_8
XFILLER_0_919 VPWR VGND sg13g2_decap_8
XFILLER_59_216 VPWR VGND sg13g2_fill_2
XFILLER_113_195 VPWR VGND sg13g2_decap_8
XFILLER_87_569 VPWR VGND sg13g2_fill_1
X_07975_ _02246_ _02248_ VPWR VGND sg13g2_inv_4
XFILLER_101_379 VPWR VGND sg13g2_decap_8
XFILLER_56_923 VPWR VGND sg13g2_fill_2
X_09645_ _03762_ _03666_ _03655_ VPWR VGND sg13g2_nand2_1
XFILLER_55_411 VPWR VGND sg13g2_decap_8
XFILLER_83_786 VPWR VGND sg13g2_decap_4
XFILLER_43_617 VPWR VGND sg13g2_decap_8
XFILLER_35_14 VPWR VGND sg13g2_decap_8
XFILLER_27_157 VPWR VGND sg13g2_decap_4
X_09576_ _03693_ net1806 acc_sum.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_82_296 VPWR VGND sg13g2_decap_8
XFILLER_71_959 VPWR VGND sg13g2_decap_4
XFILLER_70_414 VPWR VGND sg13g2_decap_8
XFILLER_42_105 VPWR VGND sg13g2_decap_8
XFILLER_24_831 VPWR VGND sg13g2_fill_1
X_08527_ _02751_ _02749_ acc_sum.op_sign_logic0.mantisa_b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_23_330 VPWR VGND sg13g2_decap_8
X_08458_ _02682_ _02690_ _02691_ VPWR VGND sg13g2_nor2_1
Xclkbuf_5_20__f_clk clknet_4_10_0_clk clknet_5_20__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_24_897 VPWR VGND sg13g2_decap_8
X_07409_ _01748_ net1889 acc\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_51_35 VPWR VGND sg13g2_decap_8
XFILLER_109_402 VPWR VGND sg13g2_decap_8
X_08389_ _02626_ _02589_ _01360_ VPWR VGND sg13g2_nor2_1
XFILLER_13_1003 VPWR VGND sg13g2_decap_8
X_10420_ _04469_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[9\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[9\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_109_435 VPWR VGND sg13g2_decap_4
XFILLER_125_928 VPWR VGND sg13g2_decap_8
XFILLER_109_468 VPWR VGND sg13g2_decap_8
X_10351_ VPWR _04401_ _04400_ VGND sg13g2_inv_1
XFILLER_124_449 VPWR VGND sg13g2_fill_2
X_13070_ _06838_ _06816_ _06820_ VPWR VGND sg13g2_nand2b_1
XFILLER_3_735 VPWR VGND sg13g2_decap_8
X_10282_ _04351_ net1830 _04210_ _04224_ net1829 VPWR VGND sg13g2_a22oi_1
X_12021_ _05870_ VPWR _00973_ VGND net1873 _05868_ sg13g2_o21ai_1
XFILLER_120_600 VPWR VGND sg13g2_decap_8
XFILLER_78_514 VPWR VGND sg13g2_decap_8
XFILLER_120_633 VPWR VGND sg13g2_decap_8
XFILLER_116_61 VPWR VGND sg13g2_decap_8
XFILLER_120_699 VPWR VGND sg13g2_decap_8
XFILLER_46_400 VPWR VGND sg13g2_decap_8
X_13972_ VPWR _00523_ net25 VGND sg13g2_inv_1
XFILLER_19_603 VPWR VGND sg13g2_fill_2
X_12923_ _06696_ _06695_ net1922 _06697_ VPWR VGND sg13g2_a21o_2
XFILLER_74_775 VPWR VGND sg13g2_fill_1
XFILLER_74_753 VPWR VGND sg13g2_fill_2
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_46_444 VPWR VGND sg13g2_fill_1
XFILLER_18_135 VPWR VGND sg13g2_decap_8
X_12854_ _06634_ _06633_ net1960 VPWR VGND sg13g2_nand2_1
XFILLER_62_948 VPWR VGND sg13g2_fill_2
XFILLER_62_937 VPWR VGND sg13g2_decap_8
XFILLER_46_488 VPWR VGND sg13g2_decap_8
XFILLER_92_75 VPWR VGND sg13g2_fill_1
X_12785_ _06568_ _06569_ _06570_ VPWR VGND sg13g2_nor2_1
X_11805_ VGND VPWR net1758 _05705_ _05706_ _05572_ sg13g2_a21oi_1
X_14524_ _00325_ VGND VPWR _01060_ fpdiv.reg_a_out\[15\] clknet_leaf_91_clk sg13g2_dfrbpq_1
XFILLER_42_683 VPWR VGND sg13g2_decap_8
XFILLER_15_875 VPWR VGND sg13g2_decap_8
X_11736_ _05640_ _05592_ _05639_ VPWR VGND sg13g2_nand2b_1
XFILLER_42_694 VPWR VGND sg13g2_fill_1
XFILLER_41_193 VPWR VGND sg13g2_fill_2
X_14455_ _00256_ VGND VPWR _00994_ fpmul.seg_reg0.q\[40\] clknet_leaf_104_clk sg13g2_dfrbpq_1
X_11667_ _05572_ _05570_ fp16_sum_pipe.reg3en.q\[0\] VPWR VGND sg13g2_nand2_2
XFILLER_30_878 VPWR VGND sg13g2_fill_1
XFILLER_127_210 VPWR VGND sg13g2_decap_8
X_14386_ _00187_ VGND VPWR net1861 fpmul.reg3en.q\[0\] clknet_leaf_17_clk sg13g2_dfrbpq_1
X_13406_ _07081_ VPWR _00800_ VGND _07032_ net1721 sg13g2_o21ai_1
XFILLER_10_580 VPWR VGND sg13g2_fill_1
X_10618_ VPWR _04631_ _04630_ VGND sg13g2_inv_1
X_11598_ _05401_ _05423_ _05503_ VPWR VGND sg13g2_nor2_1
Xplace1718 _02650_ net1718 VPWR VGND sg13g2_buf_2
Xplace1707 _02652_ net1707 VPWR VGND sg13g2_buf_2
X_13337_ _07041_ net1726 fp16_res_pipe.x2\[10\] VPWR VGND sg13g2_nand2_1
X_10549_ _04584_ VPWR _01159_ VGND net1846 _04583_ sg13g2_o21ai_1
XFILLER_127_287 VPWR VGND sg13g2_decap_8
XFILLER_109_991 VPWR VGND sg13g2_decap_8
Xplace1729 net1728 net1729 VPWR VGND sg13g2_buf_2
XFILLER_108_490 VPWR VGND sg13g2_fill_1
X_13268_ acc\[10\] net1676 _06988_ VPWR VGND sg13g2_nor2_1
XFILLER_97_823 VPWR VGND sg13g2_fill_1
X_13199_ _06934_ net1713 sipo.word\[4\] VPWR VGND sg13g2_nand2_1
X_12219_ _06065_ net1859 net1865 VPWR VGND sg13g2_nand2_1
XFILLER_123_493 VPWR VGND sg13g2_fill_2
XFILLER_111_644 VPWR VGND sg13g2_fill_1
XFILLER_96_322 VPWR VGND sg13g2_decap_8
XFILLER_69_558 VPWR VGND sg13g2_decap_8
XFILLER_111_677 VPWR VGND sg13g2_decap_8
X_07760_ VGND VPWR _01932_ _01943_ _02063_ _02062_ sg13g2_a21oi_1
XFILLER_110_187 VPWR VGND sg13g2_fill_1
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_07691_ _01999_ _01949_ acc_sub.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_53_915 VPWR VGND sg13g2_decap_8
X_09430_ VPWR _03572_ fp16_res_pipe.add_renorm0.mantisa\[0\] VGND sg13g2_inv_1
XFILLER_53_937 VPWR VGND sg13g2_decap_8
XFILLER_37_499 VPWR VGND sg13g2_fill_1
XFILLER_24_105 VPWR VGND sg13g2_decap_4
XFILLER_80_778 VPWR VGND sg13g2_fill_1
X_09361_ _03505_ _03511_ _03504_ _01274_ VPWR VGND sg13g2_nand3_1
XFILLER_17_190 VPWR VGND sg13g2_decap_8
XFILLER_24_127 VPWR VGND sg13g2_decap_8
X_08312_ _02558_ net1778 fp16_sum_pipe.op_sign_logic0.mantisa_b\[0\] VPWR VGND sg13g2_nand2_1
X_09292_ _03445_ _03369_ _03446_ VPWR VGND sg13g2_nor2_1
X_08243_ _02495_ net1638 _02494_ VPWR VGND sg13g2_nand2_1
XFILLER_21_889 VPWR VGND sg13g2_decap_8
XFILLER_119_744 VPWR VGND sg13g2_decap_8
XFILLER_118_210 VPWR VGND sg13g2_decap_8
X_08174_ _02433_ net1774 fp16_sum_pipe.op_sign_logic0.mantisa_a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_20_399 VPWR VGND sg13g2_decap_8
X_07125_ VGND VPWR _01490_ _01492_ _01489_ _01496_ sg13g2_a21oi_1
XFILLER_21_49 VPWR VGND sg13g2_decap_8
XFILLER_0_705 VPWR VGND sg13g2_decap_8
XFILLER_114_471 VPWR VGND sg13g2_decap_8
XFILLER_99_171 VPWR VGND sg13g2_decap_8
XFILLER_88_834 VPWR VGND sg13g2_decap_4
XFILLER_102_644 VPWR VGND sg13g2_decap_4
XFILLER_87_322 VPWR VGND sg13g2_decap_8
XFILLER_48_709 VPWR VGND sg13g2_fill_2
XFILLER_102_688 VPWR VGND sg13g2_fill_2
XFILLER_75_528 VPWR VGND sg13g2_fill_2
XFILLER_75_506 VPWR VGND sg13g2_decap_8
XFILLER_101_198 VPWR VGND sg13g2_decap_8
XFILLER_101_176 VPWR VGND sg13g2_decap_8
XFILLER_56_720 VPWR VGND sg13g2_fill_2
XFILLER_28_400 VPWR VGND sg13g2_decap_8
XFILLER_28_411 VPWR VGND sg13g2_fill_1
XFILLER_29_934 VPWR VGND sg13g2_decap_8
X_07958_ VPWR _02232_ _02204_ VGND sg13g2_inv_1
X_07889_ _02171_ VPWR _01399_ VGND net1891 _02091_ sg13g2_o21ai_1
XFILLER_71_701 VPWR VGND sg13g2_decap_4
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_16_606 VPWR VGND sg13g2_fill_2
X_09628_ VGND VPWR _03704_ _03714_ _03745_ _03744_ sg13g2_a21oi_1
XFILLER_55_285 VPWR VGND sg13g2_decap_8
X_09559_ _03652_ _03655_ _03675_ _03631_ _03676_ VPWR VGND sg13g2_nor4_1
X_12570_ _06386_ _06384_ _06385_ VPWR VGND sg13g2_xnor2_1
XFILLER_52_981 VPWR VGND sg13g2_fill_2
XFILLER_52_970 VPWR VGND sg13g2_decap_8
XFILLER_43_469 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_decap_8
XFILLER_23_160 VPWR VGND sg13g2_decap_8
X_11521_ _05426_ fp16_sum_pipe.add_renorm0.mantisa\[3\] fp16_sum_pipe.add_renorm0.mantisa\[2\]
+ VPWR VGND sg13g2_nand2_2
X_11452_ _05377_ VPWR _01049_ VGND net1946 _05376_ sg13g2_o21ai_1
X_14240_ _00041_ VGND VPWR _00791_ instr\[5\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_14171_ VPWR _00722_ net103 VGND sg13g2_inv_1
X_11383_ _05333_ acc_sum.exp_mant_logic0.b\[1\] _05146_ acc_sum.exp_mant_logic0.b\[0\]
+ net1654 VPWR VGND sg13g2_a22oi_1
X_10403_ _04452_ _04392_ _04453_ VPWR VGND sg13g2_nor2_1
XFILLER_125_725 VPWR VGND sg13g2_decap_8
XFILLER_124_224 VPWR VGND sg13g2_decap_8
X_13122_ _06876_ VPWR _00879_ VGND net1862 _06732_ sg13g2_o21ai_1
XFILLER_106_950 VPWR VGND sg13g2_decap_8
XFILLER_79_801 VPWR VGND sg13g2_decap_8
XFILLER_3_532 VPWR VGND sg13g2_decap_8
XFILLER_2_0 VPWR VGND sg13g2_decap_8
X_13053_ _06821_ _06817_ _06820_ VPWR VGND sg13g2_nand2_1
XFILLER_3_587 VPWR VGND sg13g2_decap_4
X_10265_ _01194_ _04334_ _04335_ VPWR VGND sg13g2_nand2_1
XFILLER_121_931 VPWR VGND sg13g2_decap_8
XFILLER_79_856 VPWR VGND sg13g2_fill_2
XFILLER_79_845 VPWR VGND sg13g2_decap_8
X_12004_ VGND VPWR _05853_ _05856_ _05858_ _05857_ sg13g2_a21oi_1
XFILLER_120_463 VPWR VGND sg13g2_fill_2
XFILLER_78_377 VPWR VGND sg13g2_fill_1
XFILLER_66_528 VPWR VGND sg13g2_decap_4
XFILLER_66_506 VPWR VGND sg13g2_fill_1
XFILLER_120_496 VPWR VGND sg13g2_decap_8
X_13955_ VPWR _00506_ net97 VGND sg13g2_inv_1
XFILLER_35_904 VPWR VGND sg13g2_decap_8
X_12906_ _06680_ _06681_ _06671_ _00900_ VPWR VGND sg13g2_nand3_1
XFILLER_74_572 VPWR VGND sg13g2_decap_8
X_13886_ VPWR _00437_ net48 VGND sg13g2_inv_1
XFILLER_19_488 VPWR VGND sg13g2_fill_2
XFILLER_19_499 VPWR VGND sg13g2_fill_2
X_12837_ _06618_ net1909 fp16_res_pipe.y\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_62_745 VPWR VGND sg13g2_fill_1
XFILLER_50_907 VPWR VGND sg13g2_fill_2
XFILLER_34_436 VPWR VGND sg13g2_fill_1
XFILLER_50_929 VPWR VGND sg13g2_decap_8
XFILLER_15_650 VPWR VGND sg13g2_decap_4
X_12768_ _00020_ _00019_ _00018_ _00017_ _06553_ VPWR VGND sg13g2_nor4_1
X_12699_ _06507_ _06459_ _06508_ VPWR VGND sg13g2_xor2_1
X_14507_ _00308_ VGND VPWR _01043_ fpdiv.reg_b_out\[14\] clknet_leaf_91_clk sg13g2_dfrbpq_2
X_14438_ _00239_ VGND VPWR _00977_ fpmul.seg_reg0.q\[23\] clknet_leaf_93_clk sg13g2_dfrbpq_1
XFILLER_7_860 VPWR VGND sg13g2_decap_8
XFILLER_115_224 VPWR VGND sg13g2_decap_8
X_14369_ _00170_ VGND VPWR _00910_ fpmul.reg_b_out\[0\] clknet_leaf_104_clk sg13g2_dfrbpq_2
XFILLER_116_758 VPWR VGND sg13g2_decap_8
X_08930_ _03117_ _03014_ _02967_ VPWR VGND sg13g2_nand2_1
X_08861_ acc_sub.seg_reg1.q\[21\] _03047_ _03042_ _03048_ VPWR VGND sg13g2_nor3_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
XFILLER_112_964 VPWR VGND sg13g2_decap_8
X_07812_ _02110_ acc_sub.exp_mant_logic0.b\[1\] net1669 acc_sub.op_sign_logic0.mantisa_b\[4\]
+ net1781 VPWR VGND sg13g2_a22oi_1
XFILLER_97_686 VPWR VGND sg13g2_fill_2
XFILLER_97_675 VPWR VGND sg13g2_decap_4
XFILLER_69_366 VPWR VGND sg13g2_fill_1
X_08792_ acc_sub.add_renorm0.mantisa\[10\] _02978_ _02979_ VPWR VGND sg13g2_nor2_2
XFILLER_96_196 VPWR VGND sg13g2_fill_1
XFILLER_96_185 VPWR VGND sg13g2_decap_4
XFILLER_85_837 VPWR VGND sg13g2_fill_1
XFILLER_84_325 VPWR VGND sg13g2_fill_1
XFILLER_57_539 VPWR VGND sg13g2_decap_8
X_07743_ VPWR _02048_ _01959_ VGND sg13g2_inv_1
X_07674_ _01982_ _01983_ _01981_ _01984_ VPWR VGND sg13g2_nand3_1
XFILLER_93_870 VPWR VGND sg13g2_decap_8
XFILLER_53_734 VPWR VGND sg13g2_fill_1
XFILLER_26_926 VPWR VGND sg13g2_decap_8
X_09413_ _03555_ _03557_ _03554_ _01268_ VPWR VGND sg13g2_nand3_1
XFILLER_16_49 VPWR VGND sg13g2_decap_8
X_09344_ _03495_ VPWR _03496_ VGND _03391_ _03494_ sg13g2_o21ai_1
X_09275_ VGND VPWR _03428_ _03424_ _03429_ _03395_ sg13g2_a21oi_1
XFILLER_119_530 VPWR VGND sg13g2_decap_8
X_08226_ _02480_ _02338_ _02472_ VPWR VGND sg13g2_nand2_1
XFILLER_5_808 VPWR VGND sg13g2_fill_1
X_08157_ _02413_ _02416_ _02412_ _02417_ VPWR VGND sg13g2_nand3_1
XFILLER_113_7 VPWR VGND sg13g2_decap_8
X_08088_ _02354_ net1639 _02325_ VPWR VGND sg13g2_nand2b_1
XFILLER_122_728 VPWR VGND sg13g2_decap_8
XFILLER_106_268 VPWR VGND sg13g2_decap_4
XFILLER_121_238 VPWR VGND sg13g2_decap_8
XFILLER_103_953 VPWR VGND sg13g2_decap_8
X_10050_ _04138_ _04109_ _04137_ VPWR VGND sg13g2_nand2_2
XFILLER_88_664 VPWR VGND sg13g2_decap_8
XFILLER_76_804 VPWR VGND sg13g2_fill_1
XFILLER_102_474 VPWR VGND sg13g2_decap_8
XFILLER_87_174 VPWR VGND sg13g2_decap_8
XFILLER_76_859 VPWR VGND sg13g2_decap_8
XFILLER_75_336 VPWR VGND sg13g2_decap_4
XFILLER_57_56 VPWR VGND sg13g2_fill_1
XFILLER_57_89 VPWR VGND sg13g2_decap_8
XFILLER_29_742 VPWR VGND sg13g2_decap_8
XFILLER_90_339 VPWR VGND sg13g2_fill_1
XFILLER_84_881 VPWR VGND sg13g2_fill_1
XFILLER_73_22 VPWR VGND sg13g2_decap_8
X_13740_ VPWR _00291_ net52 VGND sg13g2_inv_1
XFILLER_17_926 VPWR VGND sg13g2_decap_8
X_10952_ _04956_ _03586_ _04958_ VPWR VGND sg13g2_and2_1
XFILLER_113_84 VPWR VGND sg13g2_decap_8
XFILLER_83_380 VPWR VGND sg13g2_decap_4
XFILLER_28_296 VPWR VGND sg13g2_fill_1
X_13671_ VPWR _00222_ net125 VGND sg13g2_inv_1
XFILLER_32_929 VPWR VGND sg13g2_decap_8
X_10883_ _04894_ _04851_ _04817_ VPWR VGND sg13g2_nand2_1
X_12553_ _06370_ _06354_ div_result\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_40_973 VPWR VGND sg13g2_fill_2
XFILLER_40_962 VPWR VGND sg13g2_fill_1
XFILLER_40_951 VPWR VGND sg13g2_decap_8
XFILLER_24_491 VPWR VGND sg13g2_decap_4
XFILLER_89_1007 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_11_163 VPWR VGND sg13g2_decap_8
X_11504_ _05409_ fp16_sum_pipe.add_renorm0.mantisa\[2\] VPWR VGND sg13g2_inv_2
X_12484_ _06246_ _06209_ _06322_ VPWR VGND sg13g2_nor2b_1
X_14223_ _00024_ VGND VPWR _00774_ sipo.shift_reg\[4\] clknet_leaf_14_clk sg13g2_dfrbpq_1
X_11435_ _05366_ VPWR _01055_ VGND net1937 _05365_ sg13g2_o21ai_1
X_14154_ VPWR _00705_ net131 VGND sg13g2_inv_1
XFILLER_98_52 VPWR VGND sg13g2_decap_8
X_11366_ _05318_ net1761 acc_sum.op_sign_logic0.mantisa_b\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_112_216 VPWR VGND sg13g2_fill_2
X_14085_ VPWR _00636_ net89 VGND sg13g2_inv_1
X_13105_ _06863_ VPWR _00883_ VGND net1862 _06688_ sg13g2_o21ai_1
X_11297_ _05150_ _05052_ _05256_ VPWR VGND sg13g2_nor2b_2
X_10317_ _04376_ net1911 fp16_res_pipe.x2\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_4_874 VPWR VGND sg13g2_decap_8
X_13036_ _06765_ _06802_ _06804_ VPWR VGND sg13g2_nor2_1
X_10248_ _01195_ _04318_ _04319_ VPWR VGND sg13g2_nand2_1
XFILLER_113_1005 VPWR VGND sg13g2_decap_8
XFILLER_39_517 VPWR VGND sg13g2_decap_8
X_10179_ VGND VPWR net1828 _04224_ _04258_ _04257_ sg13g2_a21oi_1
XFILLER_19_241 VPWR VGND sg13g2_decap_8
XFILLER_75_881 VPWR VGND sg13g2_fill_2
X_13938_ VPWR _00489_ net25 VGND sg13g2_inv_1
XFILLER_34_200 VPWR VGND sg13g2_decap_4
XFILLER_62_564 VPWR VGND sg13g2_fill_2
XFILLER_35_789 VPWR VGND sg13g2_decap_4
X_13869_ VPWR _00420_ net14 VGND sg13g2_inv_1
X_07390_ VPWR _01735_ acc_sub.exp_mant_logic0.a\[9\] VGND sg13g2_inv_1
XFILLER_22_428 VPWR VGND sg13g2_fill_1
XFILLER_15_491 VPWR VGND sg13g2_decap_8
X_09060_ VPWR _03245_ _03189_ VGND sg13g2_inv_1
XFILLER_31_984 VPWR VGND sg13g2_decap_8
XFILLER_120_1009 VPWR VGND sg13g2_decap_4
X_08011_ _02277_ _02264_ fp16_sum_pipe.exp_mant_logic0.b\[8\] VPWR VGND sg13g2_nand2_1
X_08913_ VPWR _03100_ _03099_ VGND sg13g2_inv_1
XFILLER_112_761 VPWR VGND sg13g2_decap_8
XFILLER_98_995 VPWR VGND sg13g2_decap_8
XFILLER_97_461 VPWR VGND sg13g2_fill_2
XFILLER_97_450 VPWR VGND sg13g2_fill_1
XFILLER_58_826 VPWR VGND sg13g2_decap_8
X_08844_ VPWR _03031_ _03030_ VGND sg13g2_inv_1
XFILLER_100_923 VPWR VGND sg13g2_decap_8
XFILLER_85_623 VPWR VGND sg13g2_decap_8
XFILLER_69_185 VPWR VGND sg13g2_decap_8
XFILLER_84_122 VPWR VGND sg13g2_decap_8
X_08775_ _02963_ acc_sum.exp_mant_logic0.a\[0\] VPWR VGND sg13g2_inv_2
X_07726_ _02031_ VPWR _02032_ VGND _01745_ _02015_ sg13g2_o21ai_1
XFILLER_72_317 VPWR VGND sg13g2_decap_8
XFILLER_38_594 VPWR VGND sg13g2_fill_1
X_07657_ _01968_ net1649 net1792 VPWR VGND sg13g2_nand2_1
XFILLER_81_884 VPWR VGND sg13g2_fill_1
XFILLER_53_575 VPWR VGND sg13g2_decap_8
XFILLER_43_14 VPWR VGND sg13g2_decap_8
X_07588_ VGND VPWR net1687 _01887_ _01902_ _01901_ sg13g2_a21oi_1
XFILLER_40_247 VPWR VGND sg13g2_decap_8
X_09327_ _03479_ VPWR _03480_ VGND _03444_ _03368_ sg13g2_o21ai_1
XFILLER_22_940 VPWR VGND sg13g2_decap_8
XFILLER_126_308 VPWR VGND sg13g2_decap_8
X_09258_ VPWR _03412_ fp16_res_pipe.op_sign_logic0.mantisa_a\[1\] VGND sg13g2_inv_1
XFILLER_107_500 VPWR VGND sg13g2_decap_4
X_09189_ _03349_ acc_sum.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_inv_2
XFILLER_5_627 VPWR VGND sg13g2_decap_8
X_08209_ _02464_ _02199_ _02463_ _02465_ VPWR VGND _02194_ sg13g2_nand4_1
X_11220_ _05179_ _05184_ _05185_ _05186_ VPWR VGND sg13g2_nor3_1
XFILLER_49_1013 VPWR VGND sg13g2_fill_1
XFILLER_49_1002 VPWR VGND sg13g2_decap_8
XFILLER_4_126 VPWR VGND sg13g2_decap_8
X_11151_ _05116_ _05120_ _05121_ VPWR VGND sg13g2_nor2_1
XFILLER_89_951 VPWR VGND sg13g2_decap_8
Xplace1890 net1889 net1890 VPWR VGND sg13g2_buf_1
XFILLER_1_822 VPWR VGND sg13g2_decap_8
X_10102_ _03611_ _04124_ _04186_ VPWR VGND sg13g2_nor2_1
XFILLER_103_761 VPWR VGND sg13g2_decap_8
X_11082_ _05058_ _05052_ acc_sum.exp_mant_logic0.a\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_49_815 VPWR VGND sg13g2_fill_1
X_14910_ _00711_ VGND VPWR _01430_ acc_sub.op_sign_logic0.mantisa_a\[9\] clknet_leaf_62_clk
+ sg13g2_dfrbpq_1
XFILLER_103_783 VPWR VGND sg13g2_fill_2
XFILLER_49_826 VPWR VGND sg13g2_decap_8
XFILLER_0_365 VPWR VGND sg13g2_decap_8
XFILLER_1_899 VPWR VGND sg13g2_decap_8
X_10033_ _04115_ _04120_ _04121_ VPWR VGND sg13g2_nor2_1
XFILLER_102_282 VPWR VGND sg13g2_decap_4
XFILLER_64_807 VPWR VGND sg13g2_fill_2
X_14841_ _00642_ VGND VPWR _01365_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[3\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
XFILLER_84_43 VPWR VGND sg13g2_fill_1
XFILLER_75_188 VPWR VGND sg13g2_fill_2
XFILLER_1_1004 VPWR VGND sg13g2_decap_8
X_14772_ _00573_ VGND VPWR _01296_ acc_sub.y\[1\] clknet_leaf_46_clk sg13g2_dfrbpq_1
X_11984_ fpmul.reg_b_out\[9\] fpmul.reg_a_out\[9\] _05838_ VPWR VGND sg13g2_xor2_1
XFILLER_16_222 VPWR VGND sg13g2_decap_8
XFILLER_29_594 VPWR VGND sg13g2_fill_1
X_13723_ VPWR _00274_ net139 VGND sg13g2_inv_1
XFILLER_16_255 VPWR VGND sg13g2_fill_1
XFILLER_16_266 VPWR VGND sg13g2_decap_8
XFILLER_17_70 VPWR VGND sg13g2_decap_8
XFILLER_17_81 VPWR VGND sg13g2_fill_1
X_10935_ _04942_ _04941_ _04846_ VPWR VGND sg13g2_nand2b_1
X_13654_ VPWR _00205_ net70 VGND sg13g2_inv_1
XFILLER_16_299 VPWR VGND sg13g2_decap_8
X_10866_ _04878_ _04875_ _04877_ VPWR VGND sg13g2_nand2_1
X_12605_ net1851 _06421_ VPWR VGND sg13g2_inv_4
XFILLER_13_940 VPWR VGND sg13g2_decap_8
X_13585_ VPWR _00136_ net115 VGND sg13g2_inv_1
X_10797_ _04809_ _04808_ VPWR VGND sg13g2_inv_2
XFILLER_117_308 VPWR VGND sg13g2_fill_2
XFILLER_40_792 VPWR VGND sg13g2_fill_2
XFILLER_8_432 VPWR VGND sg13g2_decap_8
XFILLER_9_955 VPWR VGND sg13g2_decap_8
XFILLER_12_483 VPWR VGND sg13g2_decap_8
XFILLER_126_820 VPWR VGND sg13g2_decap_8
X_12467_ _06309_ _06308_ _06020_ VPWR VGND sg13g2_nand2_1
XFILLER_8_476 VPWR VGND sg13g2_decap_8
X_14206_ VPWR _00757_ net132 VGND sg13g2_inv_1
X_11418_ _05355_ VPWR _01061_ VGND _05353_ fpdiv.divider0.en_r sg13g2_o21ai_1
XFILLER_126_897 VPWR VGND sg13g2_decap_8
XFILLER_99_715 VPWR VGND sg13g2_decap_8
X_14137_ VPWR _00688_ net114 VGND sg13g2_inv_1
X_12398_ _06244_ _06243_ _06207_ VPWR VGND sg13g2_nand2_1
XFILLER_4_671 VPWR VGND sg13g2_decap_8
XFILLER_98_225 VPWR VGND sg13g2_decap_8
X_11349_ _05302_ _05181_ net1812 VPWR VGND sg13g2_nand2_1
X_14068_ VPWR _00619_ net95 VGND sg13g2_inv_1
XFILLER_121_580 VPWR VGND sg13g2_fill_1
XFILLER_95_932 VPWR VGND sg13g2_decap_8
X_13019_ VPWR _06787_ _06786_ VGND sg13g2_inv_1
XFILLER_66_144 VPWR VGND sg13g2_decap_8
XFILLER_94_475 VPWR VGND sg13g2_decap_8
XFILLER_82_604 VPWR VGND sg13g2_decap_8
XFILLER_48_870 VPWR VGND sg13g2_decap_8
XFILLER_39_369 VPWR VGND sg13g2_fill_2
X_08560_ VGND VPWR _02783_ _02778_ _02784_ _02777_ sg13g2_a21oi_1
XFILLER_81_147 VPWR VGND sg13g2_fill_1
XFILLER_63_840 VPWR VGND sg13g2_decap_8
XFILLER_54_339 VPWR VGND sg13g2_fill_2
X_08491_ _02718_ VPWR _01351_ VGND net1705 _02717_ sg13g2_o21ai_1
X_07511_ _01833_ _01832_ _01802_ VPWR VGND sg13g2_nand2_1
XFILLER_81_158 VPWR VGND sg13g2_decap_8
XFILLER_35_575 VPWR VGND sg13g2_decap_8
X_07442_ _01771_ VPWR _01446_ VGND _01770_ net1750 sg13g2_o21ai_1
XFILLER_62_394 VPWR VGND sg13g2_decap_8
XFILLER_50_534 VPWR VGND sg13g2_decap_8
Xfanout18 net24 net18 VPWR VGND sg13g2_buf_1
Xfanout29 net30 net29 VPWR VGND sg13g2_buf_2
XFILLER_35_597 VPWR VGND sg13g2_decap_4
Xclkbuf_5_1__f_clk clknet_4_0_0_clk clknet_5_1__leaf_clk VPWR VGND sg13g2_buf_8
X_07373_ acc_sub.exp_mant_logic0.a\[15\] net1893 _01724_ VPWR VGND sg13g2_nor2_1
X_09112_ _03293_ VPWR _01305_ VGND net1801 _03283_ sg13g2_o21ai_1
XFILLER_13_28 VPWR VGND sg13g2_decap_8
XFILLER_31_781 VPWR VGND sg13g2_decap_4
X_09043_ _03223_ _03228_ _03229_ VPWR VGND sg13g2_nor2_1
XFILLER_117_886 VPWR VGND sg13g2_decap_8
XFILLER_116_352 VPWR VGND sg13g2_decap_8
XFILLER_2_608 VPWR VGND sg13g2_decap_8
XFILLER_86_910 VPWR VGND sg13g2_decap_8
X_09945_ VPWR _04041_ _04004_ VGND sg13g2_inv_1
X_09876_ acc_sum.y\[3\] _03757_ net1820 _01228_ VPWR VGND sg13g2_mux2_1
XFILLER_38_14 VPWR VGND sg13g2_decap_8
X_08827_ _02995_ _03013_ _03009_ _03014_ VPWR VGND sg13g2_nor3_2
XFILLER_86_987 VPWR VGND sg13g2_decap_8
XFILLER_72_103 VPWR VGND sg13g2_fill_1
XFILLER_58_689 VPWR VGND sg13g2_fill_2
XFILLER_57_155 VPWR VGND sg13g2_fill_2
XFILLER_46_829 VPWR VGND sg13g2_decap_8
X_08758_ _02952_ acc\[6\] net1896 VPWR VGND sg13g2_nand2_1
X_07709_ _01743_ _02015_ _02016_ VPWR VGND sg13g2_nor2_1
X_08689_ _02904_ _02902_ _02903_ _02823_ net1739 VPWR VGND sg13g2_a22oi_1
XFILLER_54_862 VPWR VGND sg13g2_decap_8
XFILLER_54_35 VPWR VGND sg13g2_decap_8
XFILLER_81_670 VPWR VGND sg13g2_decap_4
XFILLER_53_372 VPWR VGND sg13g2_fill_2
XFILLER_53_361 VPWR VGND sg13g2_decap_8
X_10720_ _04686_ _04702_ _04708_ _04732_ _04733_ VPWR VGND sg13g2_nor4_1
XFILLER_13_258 VPWR VGND sg13g2_decap_8
XFILLER_16_1001 VPWR VGND sg13g2_decap_8
XFILLER_110_63 VPWR VGND sg13g2_decap_8
X_10651_ _04664_ _04662_ VPWR VGND sg13g2_inv_2
XFILLER_16_1012 VPWR VGND sg13g2_fill_2
XFILLER_70_45 VPWR VGND sg13g2_decap_4
X_13370_ _07061_ net1694 sipo.word\[13\] VPWR VGND sg13g2_nand2_1
X_10582_ _04604_ acc_sub.x2\[8\] net1926 VPWR VGND sg13g2_nand2_1
XFILLER_10_954 VPWR VGND sg13g2_decap_8
XFILLER_126_105 VPWR VGND sg13g2_decap_8
X_12321_ VGND VPWR _06166_ _06167_ _06164_ _06162_ sg13g2_a21oi_2
X_12252_ _06098_ _06096_ _06097_ VPWR VGND sg13g2_nand2_1
XFILLER_6_969 VPWR VGND sg13g2_decap_8
XFILLER_108_864 VPWR VGND sg13g2_fill_1
XFILLER_102_0 VPWR VGND sg13g2_decap_8
X_11203_ _05168_ _05169_ _05167_ _05170_ VPWR VGND sg13g2_nand3_1
XFILLER_5_457 VPWR VGND sg13g2_decap_8
XFILLER_123_834 VPWR VGND sg13g2_decap_8
X_12183_ _06029_ fpmul.reg_a_out\[6\] net1864 VPWR VGND sg13g2_nand2_1
XFILLER_95_206 VPWR VGND sg13g2_fill_2
X_11134_ _05103_ _05010_ _05104_ VPWR VGND sg13g2_xor2_1
XFILLER_110_517 VPWR VGND sg13g2_decap_8
XFILLER_89_781 VPWR VGND sg13g2_fill_2
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_77_976 VPWR VGND sg13g2_decap_4
XFILLER_37_807 VPWR VGND sg13g2_decap_8
X_10016_ _04104_ _04097_ _04103_ VPWR VGND sg13g2_nand2_1
XFILLER_95_97 VPWR VGND sg13g2_fill_2
X_14824_ _00625_ VGND VPWR _01348_ acc_sum.seg_reg1.q\[21\] clknet_leaf_34_clk sg13g2_dfrbpq_1
XFILLER_92_946 VPWR VGND sg13g2_decap_8
XFILLER_28_91 VPWR VGND sg13g2_decap_4
XFILLER_91_478 VPWR VGND sg13g2_decap_4
X_14755_ _00556_ VGND VPWR _01279_ acc_sum.exp_mant_logic0.b\[0\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
X_11967_ _05822_ net1884 fpmul.reg_b_out\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_60_821 VPWR VGND sg13g2_decap_8
X_13706_ VPWR _00257_ net63 VGND sg13g2_inv_1
X_10918_ _04897_ _04926_ _04923_ _04927_ VPWR VGND sg13g2_nand3_1
XFILLER_60_854 VPWR VGND sg13g2_decap_8
X_11898_ VPWR _05779_ fpmul.seg_reg0.q\[50\] VGND sg13g2_inv_1
X_14686_ _00487_ VGND VPWR _01214_ fp16_res_pipe.seg_reg0.q\[23\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_1
XFILLER_32_556 VPWR VGND sg13g2_decap_8
X_13637_ VPWR _00188_ net124 VGND sg13g2_inv_1
X_10849_ net1825 _03580_ _04861_ VPWR VGND sg13g2_nor2_1
X_13568_ VPWR _00119_ net33 VGND sg13g2_inv_1
XFILLER_117_105 VPWR VGND sg13g2_decap_8
X_12519_ fpmul.reg_a_out\[7\] net1951 _06345_ VPWR VGND sg13g2_nor2_1
X_13499_ VPWR _00050_ net37 VGND sg13g2_inv_1
XFILLER_125_182 VPWR VGND sg13g2_decap_8
XFILLER_114_867 VPWR VGND sg13g2_decap_8
X_07991_ _02258_ VPWR _01384_ VGND _02216_ _02248_ sg13g2_o21ai_1
XFILLER_5_84 VPWR VGND sg13g2_decap_8
XFILLER_4_490 VPWR VGND sg13g2_decap_8
X_09730_ _03846_ _03840_ _03842_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_4_7_0_clk clknet_0_clk clknet_4_7_0_clk VPWR VGND sg13g2_buf_8
XFILLER_68_965 VPWR VGND sg13g2_decap_8
XFILLER_39_133 VPWR VGND sg13g2_decap_8
X_09661_ _03740_ _03777_ _03778_ VPWR VGND sg13g2_nor2_1
XFILLER_95_773 VPWR VGND sg13g2_fill_2
XFILLER_95_762 VPWR VGND sg13g2_decap_8
XFILLER_82_401 VPWR VGND sg13g2_decap_8
XFILLER_28_829 VPWR VGND sg13g2_fill_2
X_09592_ VGND VPWR net1805 _03673_ _03709_ _03708_ sg13g2_a21oi_1
XFILLER_94_294 VPWR VGND sg13g2_fill_1
X_08612_ _02835_ _02834_ _02791_ VPWR VGND sg13g2_nand2_1
XFILLER_83_946 VPWR VGND sg13g2_decap_8
XFILLER_54_103 VPWR VGND sg13g2_decap_4
X_08543_ VPWR _02767_ _02766_ VGND sg13g2_inv_1
XFILLER_54_158 VPWR VGND sg13g2_decap_8
XFILLER_39_1012 VPWR VGND sg13g2_fill_2
X_08474_ _02705_ fpdiv.divider0.remainder_reg\[9\] net1708 _01756_ fpdiv.divider0.dividend\[9\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_51_865 VPWR VGND sg13g2_decap_8
XFILLER_23_556 VPWR VGND sg13g2_decap_8
XFILLER_24_49 VPWR VGND sg13g2_decap_8
X_07425_ _01451_ _01758_ _01759_ VPWR VGND sg13g2_nand2_1
X_07356_ _01713_ acc_sub.add_renorm0.exp\[5\] VPWR VGND sg13g2_inv_2
X_07287_ _01654_ VPWR _01655_ VGND _01636_ _01650_ sg13g2_o21ai_1
X_09026_ _03097_ VPWR _03212_ VGND _03193_ _03211_ sg13g2_o21ai_1
XFILLER_3_917 VPWR VGND sg13g2_decap_8
XFILLER_123_119 VPWR VGND sg13g2_decap_8
XFILLER_117_694 VPWR VGND sg13g2_fill_2
XFILLER_104_322 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_2_416 VPWR VGND sg13g2_decap_8
XFILLER_104_355 VPWR VGND sg13g2_decap_4
XFILLER_78_707 VPWR VGND sg13g2_fill_1
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_120_848 VPWR VGND sg13g2_decap_8
X_09928_ _04025_ _04023_ _04024_ VPWR VGND sg13g2_nand2_1
X_09859_ VGND VPWR _03665_ _03844_ _03968_ _03740_ sg13g2_a21oi_1
XFILLER_85_250 VPWR VGND sg13g2_decap_8
XFILLER_74_924 VPWR VGND sg13g2_decap_8
XFILLER_46_604 VPWR VGND sg13g2_decap_8
XFILLER_105_96 VPWR VGND sg13g2_decap_8
X_12870_ _06647_ _06648_ _06638_ _00903_ VPWR VGND sg13g2_nand3_1
XFILLER_65_56 VPWR VGND sg13g2_fill_2
XFILLER_45_147 VPWR VGND sg13g2_decap_8
X_11821_ VGND VPWR _05720_ _05633_ _05721_ _05592_ sg13g2_a21oi_1
XFILLER_73_489 VPWR VGND sg13g2_fill_2
X_14540_ _00341_ VGND VPWR _01076_ acc_sum.op_sign_logic0.mantisa_b\[3\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
XFILLER_42_810 VPWR VGND sg13g2_decap_8
XFILLER_14_512 VPWR VGND sg13g2_decap_4
XFILLER_121_84 VPWR VGND sg13g2_decap_8
XFILLER_42_843 VPWR VGND sg13g2_decap_8
X_11752_ VGND VPWR _05602_ net1839 _05656_ _05655_ sg13g2_a21oi_1
XFILLER_14_545 VPWR VGND sg13g2_decap_4
X_14471_ _00272_ VGND VPWR _01010_ fpdiv.divider0.counter\[1\] clknet_leaf_73_clk
+ sg13g2_dfrbpq_1
XFILLER_81_77 VPWR VGND sg13g2_fill_1
XFILLER_41_364 VPWR VGND sg13g2_decap_8
X_11683_ net1727 _05582_ _05586_ _05587_ VPWR VGND sg13g2_a21o_2
X_10703_ _04711_ _04714_ _04716_ VPWR VGND _04627_ sg13g2_nand3b_1
X_13422_ _07090_ net1719 instr\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_41_397 VPWR VGND sg13g2_decap_8
XFILLER_41_386 VPWR VGND sg13g2_fill_1
X_10634_ _04647_ _04644_ _04646_ VPWR VGND sg13g2_xnor2_1
X_13353_ _07050_ VPWR _00822_ VGND _07006_ net1723 sg13g2_o21ai_1
XFILLER_14_82 VPWR VGND sg13g2_fill_2
XFILLER_127_458 VPWR VGND sg13g2_decap_8
X_12304_ VPWR _06150_ _06114_ VGND sg13g2_inv_1
X_10565_ VPWR _04595_ fp16_sum_pipe.add_renorm0.exp\[0\] VGND sg13g2_inv_1
XFILLER_127_469 VPWR VGND sg13g2_fill_1
XFILLER_108_661 VPWR VGND sg13g2_decap_8
X_13284_ _06999_ _06952_ _07000_ VPWR VGND sg13g2_nor2_1
XFILLER_5_254 VPWR VGND sg13g2_fill_2
X_10496_ VPWR _04541_ _04492_ VGND sg13g2_inv_1
XFILLER_114_119 VPWR VGND sg13g2_decap_8
XFILLER_107_160 VPWR VGND sg13g2_fill_2
X_12235_ _06073_ _06080_ _06081_ VPWR VGND sg13g2_nor2_1
XFILLER_30_70 VPWR VGND sg13g2_decap_8
X_12166_ _06012_ _06009_ _06010_ VPWR VGND sg13g2_nand2_1
XFILLER_2_961 VPWR VGND sg13g2_decap_8
XFILLER_68_217 VPWR VGND sg13g2_decap_8
X_11117_ VPWR _05087_ _05086_ VGND sg13g2_inv_1
XFILLER_39_7 VPWR VGND sg13g2_decap_8
XFILLER_1_471 VPWR VGND sg13g2_decap_8
XFILLER_122_196 VPWR VGND sg13g2_decap_8
XFILLER_111_859 VPWR VGND sg13g2_decap_8
XFILLER_77_751 VPWR VGND sg13g2_decap_8
X_12097_ _05943_ _05942_ _05898_ VPWR VGND sg13g2_nand2_1
XFILLER_49_464 VPWR VGND sg13g2_decap_8
X_14807_ _00608_ VGND VPWR _01331_ acc_sum.add_renorm0.exp\[4\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_80_916 VPWR VGND sg13g2_decap_8
XFILLER_91_275 VPWR VGND sg13g2_fill_1
XFILLER_91_264 VPWR VGND sg13g2_decap_8
X_12999_ _06767_ net1755 fpmul.seg_reg0.q\[13\] VPWR VGND sg13g2_nand2b_1
XFILLER_64_489 VPWR VGND sg13g2_fill_1
X_14738_ _00539_ VGND VPWR _01266_ fp16_res_pipe.add_renorm0.mantisa\[1\] clknet_leaf_136_clk
+ sg13g2_dfrbpq_1
XFILLER_17_394 VPWR VGND sg13g2_fill_1
X_14669_ _00470_ VGND VPWR _01197_ fp16_res_pipe.op_sign_logic0.mantisa_b\[6\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_2
XFILLER_32_342 VPWR VGND sg13g2_decap_8
X_07210_ _01582_ _01551_ _01549_ VPWR VGND sg13g2_nand2_2
X_08190_ _02268_ _02396_ _02447_ VPWR VGND sg13g2_nor2_1
XFILLER_119_926 VPWR VGND sg13g2_decap_8
X_07141_ _01510_ _01512_ _01513_ VPWR VGND sg13g2_nor2_2
XFILLER_118_447 VPWR VGND sg13g2_decap_8
XFILLER_69_1005 VPWR VGND sg13g2_decap_8
XFILLER_65_0 VPWR VGND sg13g2_decap_8
XFILLER_127_981 VPWR VGND sg13g2_decap_8
XFILLER_99_353 VPWR VGND sg13g2_decap_8
XFILLER_87_537 VPWR VGND sg13g2_fill_1
XFILLER_87_526 VPWR VGND sg13g2_decap_8
XFILLER_87_548 VPWR VGND sg13g2_decap_8
XFILLER_83_710 VPWR VGND sg13g2_fill_1
XFILLER_74_209 VPWR VGND sg13g2_decap_8
XFILLER_19_49 VPWR VGND sg13g2_decap_8
XFILLER_110_892 VPWR VGND sg13g2_decap_8
X_09644_ _03761_ _03630_ _03652_ VPWR VGND sg13g2_nand2_1
XFILLER_82_242 VPWR VGND sg13g2_decap_8
XFILLER_71_916 VPWR VGND sg13g2_decap_8
XFILLER_56_968 VPWR VGND sg13g2_fill_1
X_09575_ VPWR _03692_ _03691_ VGND sg13g2_inv_1
XFILLER_82_264 VPWR VGND sg13g2_fill_1
XFILLER_55_489 VPWR VGND sg13g2_fill_1
X_08526_ acc_sum.op_sign_logic0.mantisa_b\[3\] _02749_ _02750_ VPWR VGND sg13g2_nor2_1
X_08457_ fpdiv.divider0.remainder_reg\[11\] _02681_ _02690_ VPWR VGND sg13g2_nor2_1
X_07408_ _01747_ acc_sub.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_inv_2
XFILLER_51_14 VPWR VGND sg13g2_decap_8
XFILLER_50_161 VPWR VGND sg13g2_decap_8
XFILLER_11_537 VPWR VGND sg13g2_decap_8
XFILLER_23_386 VPWR VGND sg13g2_fill_1
X_08388_ VGND VPWR _02618_ _02563_ _02626_ _02625_ sg13g2_a21oi_1
XFILLER_11_559 VPWR VGND sg13g2_decap_8
X_07339_ VPWR _01700_ acc_sub.add_renorm0.mantisa\[1\] VGND sg13g2_inv_1
XFILLER_100_1007 VPWR VGND sg13g2_decap_8
XFILLER_125_907 VPWR VGND sg13g2_decap_8
X_10350_ _04400_ _04398_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[7\] VPWR VGND sg13g2_nand2_1
X_09009_ VPWR _03195_ _03187_ VGND sg13g2_inv_1
XFILLER_118_992 VPWR VGND sg13g2_decap_8
X_10281_ _04349_ VPWR _04350_ VGND _04300_ _04227_ sg13g2_o21ai_1
XFILLER_105_664 VPWR VGND sg13g2_decap_4
XFILLER_105_653 VPWR VGND sg13g2_fill_2
X_12020_ net1875 _05869_ _05870_ VPWR VGND _05846_ sg13g2_nand3b_1
XFILLER_116_40 VPWR VGND sg13g2_decap_8
XFILLER_105_686 VPWR VGND sg13g2_decap_8
XFILLER_2_279 VPWR VGND sg13g2_decap_8
XFILLER_120_645 VPWR VGND sg13g2_fill_1
XFILLER_59_784 VPWR VGND sg13g2_decap_8
XFILLER_59_773 VPWR VGND sg13g2_decap_8
XFILLER_59_762 VPWR VGND sg13g2_fill_2
XFILLER_47_924 VPWR VGND sg13g2_decap_8
X_13971_ VPWR _00522_ net25 VGND sg13g2_inv_1
XFILLER_101_892 VPWR VGND sg13g2_decap_8
XFILLER_86_581 VPWR VGND sg13g2_decap_8
XFILLER_74_710 VPWR VGND sg13g2_fill_1
X_12922_ _06696_ fp16_res_pipe.reg1en.d\[0\] fp16_res_pipe.y\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_19_648 VPWR VGND sg13g2_decap_8
XFILLER_92_21 VPWR VGND sg13g2_decap_4
XFILLER_73_231 VPWR VGND sg13g2_fill_1
XFILLER_62_905 VPWR VGND sg13g2_fill_2
XFILLER_19_659 VPWR VGND sg13g2_fill_2
XFILLER_92_43 VPWR VGND sg13g2_decap_8
X_12853_ VPWR _06633_ fpmul.reg_p_out\[10\] VGND sg13g2_inv_1
XFILLER_55_990 VPWR VGND sg13g2_fill_2
XFILLER_33_106 VPWR VGND sg13g2_decap_8
X_12784_ _06569_ piso.tx_bit_counter\[1\] piso.tx_bit_counter\[0\] VPWR VGND sg13g2_nand2_1
X_11804_ _05705_ _05704_ _05669_ VPWR VGND sg13g2_nand2b_1
XFILLER_14_320 VPWR VGND sg13g2_decap_4
XFILLER_14_331 VPWR VGND sg13g2_fill_2
XFILLER_15_854 VPWR VGND sg13g2_decap_8
XFILLER_26_180 VPWR VGND sg13g2_decap_4
XFILLER_70_982 VPWR VGND sg13g2_fill_1
X_14523_ _00324_ VGND VPWR _01059_ fpdiv.reg_a_out\[14\] clknet_leaf_91_clk sg13g2_dfrbpq_2
X_11735_ _05639_ _05596_ _05632_ VPWR VGND sg13g2_xnor2_1
X_14454_ _00255_ VGND VPWR _00993_ fpmul.seg_reg0.q\[39\] clknet_leaf_104_clk sg13g2_dfrbpq_1
X_13405_ _07081_ net1721 instr\[14\] VPWR VGND sg13g2_nand2_1
X_14385_ _00186_ VGND VPWR net1873 fpmul.reg2en.q\[0\] clknet_leaf_95_clk sg13g2_dfrbpq_2
X_10617_ VGND VPWR net1823 _04628_ _04630_ _04629_ sg13g2_a21oi_1
X_11597_ _05501_ VPWR _05502_ VGND fp16_sum_pipe.add_renorm0.mantisa\[11\] _05436_
+ sg13g2_o21ai_1
XFILLER_127_266 VPWR VGND sg13g2_decap_8
XFILLER_109_970 VPWR VGND sg13g2_decap_8
Xplace1708 _02652_ net1708 VPWR VGND sg13g2_buf_2
X_13336_ VPWR _07040_ sipo.word\[10\] VGND sg13g2_inv_1
XFILLER_41_91 VPWR VGND sg13g2_decap_8
XFILLER_6_530 VPWR VGND sg13g2_decap_8
X_10548_ _04584_ fp16_sum_pipe.seg_reg0.q\[28\] net1845 VPWR VGND sg13g2_nand2_1
XFILLER_115_428 VPWR VGND sg13g2_fill_2
XFILLER_108_480 VPWR VGND sg13g2_fill_2
X_13267_ VPWR VGND acc_sum.y\[10\] _06986_ net1729 net1743 _06987_ sipo.word\[10\]
+ sg13g2_a221oi_1
Xplace1719 _07076_ net1719 VPWR VGND sg13g2_buf_2
XFILLER_97_802 VPWR VGND sg13g2_decap_8
X_12218_ _06064_ net1858 net1866 VPWR VGND sg13g2_nand2_1
X_10479_ VGND VPWR net1673 _04523_ _04526_ _04525_ sg13g2_a21oi_1
XFILLER_29_1011 VPWR VGND sg13g2_fill_2
XFILLER_124_984 VPWR VGND sg13g2_decap_8
XFILLER_116_1003 VPWR VGND sg13g2_decap_8
X_13198_ VPWR _06933_ sipo.shift_reg\[5\] VGND sg13g2_inv_1
XFILLER_111_656 VPWR VGND sg13g2_decap_8
X_12149_ _05995_ net1855 net1864 VPWR VGND sg13g2_nand2_1
XFILLER_110_133 VPWR VGND sg13g2_fill_1
XFILLER_84_529 VPWR VGND sg13g2_fill_1
XFILLER_77_581 VPWR VGND sg13g2_decap_8
XFILLER_49_272 VPWR VGND sg13g2_decap_8
XFILLER_37_401 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_07690_ _01425_ _01997_ _01998_ VPWR VGND sg13g2_nand2_1
XFILLER_53_905 VPWR VGND sg13g2_decap_8
XFILLER_37_445 VPWR VGND sg13g2_decap_8
XFILLER_92_595 VPWR VGND sg13g2_decap_8
XFILLER_80_713 VPWR VGND sg13g2_decap_4
XFILLER_52_415 VPWR VGND sg13g2_decap_8
X_09360_ _03511_ _03510_ _03501_ VPWR VGND sg13g2_nand2_1
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
X_08311_ _02557_ net1638 _02556_ VPWR VGND sg13g2_nand2_1
X_09291_ fp16_res_pipe.op_sign_logic0.mantisa_b\[10\] _03444_ _03445_ VPWR VGND sg13g2_nor2_1
X_08242_ _02492_ _02493_ _02491_ _02494_ VPWR VGND sg13g2_nand3_1
XFILLER_21_846 VPWR VGND sg13g2_decap_8
XFILLER_32_161 VPWR VGND sg13g2_fill_2
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_119_723 VPWR VGND sg13g2_decap_8
XFILLER_32_194 VPWR VGND sg13g2_decap_8
X_08173_ _02432_ _02431_ net1639 VPWR VGND sg13g2_nand2_1
XFILLER_20_378 VPWR VGND sg13g2_fill_2
XFILLER_21_28 VPWR VGND sg13g2_decap_8
XFILLER_118_266 VPWR VGND sg13g2_decap_8
XFILLER_107_929 VPWR VGND sg13g2_decap_8
XFILLER_118_277 VPWR VGND sg13g2_fill_2
XFILLER_115_984 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_87_345 VPWR VGND sg13g2_fill_1
XFILLER_101_144 VPWR VGND sg13g2_decap_8
XFILLER_29_913 VPWR VGND sg13g2_decap_8
X_07957_ VGND VPWR _02229_ _02230_ _02231_ _02209_ sg13g2_a21oi_1
XFILLER_87_389 VPWR VGND sg13g2_fill_1
XFILLER_46_14 VPWR VGND sg13g2_decap_8
X_07888_ _02171_ net1891 acc_sub.x2\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_83_551 VPWR VGND sg13g2_decap_8
X_09627_ VGND VPWR _03704_ _03710_ _03744_ _03714_ sg13g2_a21oi_1
XFILLER_83_595 VPWR VGND sg13g2_decap_8
XFILLER_83_562 VPWR VGND sg13g2_fill_2
XFILLER_70_201 VPWR VGND sg13g2_decap_8
XFILLER_44_949 VPWR VGND sg13g2_decap_4
XFILLER_16_629 VPWR VGND sg13g2_fill_1
XFILLER_28_489 VPWR VGND sg13g2_decap_4
X_09558_ VPWR _03675_ _03674_ VGND sg13g2_inv_1
XFILLER_70_245 VPWR VGND sg13g2_fill_2
XFILLER_70_234 VPWR VGND sg13g2_decap_8
XFILLER_70_212 VPWR VGND sg13g2_fill_2
XFILLER_102_97 VPWR VGND sg13g2_decap_4
X_08509_ acc_sum.op_sign_logic0.mantisa_a\[8\] acc_sum.op_sign_logic0.mantisa_b\[8\]
+ _02733_ VPWR VGND sg13g2_nor2b_2
XFILLER_24_640 VPWR VGND sg13g2_fill_2
XFILLER_11_301 VPWR VGND sg13g2_decap_4
X_11520_ VPWR _05425_ fp16_sum_pipe.add_renorm0.mantisa\[4\] VGND sg13g2_inv_1
X_09489_ _03610_ VPWR _01245_ VGND net1918 _03609_ sg13g2_o21ai_1
XFILLER_7_305 VPWR VGND sg13g2_fill_2
XFILLER_11_356 VPWR VGND sg13g2_decap_8
X_11451_ _05377_ acc_sub.x2\[4\] net1946 VPWR VGND sg13g2_nand2_1
XFILLER_8_839 VPWR VGND sg13g2_decap_8
XFILLER_11_367 VPWR VGND sg13g2_fill_2
X_14170_ VPWR _00721_ net132 VGND sg13g2_inv_1
X_11382_ _05332_ acc_sum.exp_mant_logic0.b\[3\] _05192_ acc_sum.exp_mant_logic0.b\[2\]
+ _05181_ VPWR VGND sg13g2_a22oi_1
X_10402_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[8\] _04390_ _04452_ VPWR VGND sg13g2_nor2_1
XFILLER_124_203 VPWR VGND sg13g2_decap_8
X_13121_ net1700 _06875_ _06802_ _06876_ VPWR VGND sg13g2_nand3_1
XFILLER_3_511 VPWR VGND sg13g2_decap_8
X_10333_ fp16_sum_pipe.op_sign_logic0.s_b fp16_sum_pipe.op_sign_logic0.s_a _04384_
+ VPWR VGND sg13g2_xor2_1
XFILLER_121_910 VPWR VGND sg13g2_decap_8
XFILLER_105_472 VPWR VGND sg13g2_decap_8
XFILLER_87_21 VPWR VGND sg13g2_fill_1
X_13052_ _06819_ fpmul.seg_reg0.q\[23\] _06820_ VPWR VGND sg13g2_xor2_1
X_10264_ _04335_ fp16_res_pipe.exp_mant_logic0.b\[0\] net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[3\]
+ _03988_ VPWR VGND sg13g2_a22oi_1
X_12003_ _05854_ _05855_ _05857_ VPWR VGND sg13g2_nor2b_1
X_10195_ _04149_ _04056_ _04272_ VPWR VGND sg13g2_nor2b_1
XFILLER_121_987 VPWR VGND sg13g2_decap_8
XFILLER_94_816 VPWR VGND sg13g2_decap_4
XFILLER_87_98 VPWR VGND sg13g2_decap_8
XFILLER_78_389 VPWR VGND sg13g2_fill_1
X_13954_ VPWR _00505_ net79 VGND sg13g2_inv_1
XFILLER_47_765 VPWR VGND sg13g2_fill_2
X_12905_ _06681_ net1717 _00011_ VPWR VGND sg13g2_nand2_1
XFILLER_46_253 VPWR VGND sg13g2_decap_8
X_13885_ VPWR _00436_ net48 VGND sg13g2_inv_1
XFILLER_19_467 VPWR VGND sg13g2_decap_8
X_12836_ acc\[11\] net1908 net1767 _06617_ VPWR VGND sg13g2_nand3_1
XFILLER_36_91 VPWR VGND sg13g2_decap_8
XFILLER_34_459 VPWR VGND sg13g2_decap_8
XFILLER_34_426 VPWR VGND sg13g2_decap_4
XFILLER_62_779 VPWR VGND sg13g2_decap_4
XFILLER_61_245 VPWR VGND sg13g2_decap_8
XFILLER_43_971 VPWR VGND sg13g2_decap_4
X_12767_ _00016_ _00015_ _00014_ _00013_ _06552_ VPWR VGND sg13g2_nor4_1
XFILLER_70_790 VPWR VGND sg13g2_fill_1
X_14506_ _00307_ VGND VPWR _01042_ fpdiv.reg_b_out\[13\] clknet_leaf_91_clk sg13g2_dfrbpq_1
XFILLER_15_695 VPWR VGND sg13g2_decap_8
XFILLER_30_621 VPWR VGND sg13g2_decap_8
XFILLER_30_632 VPWR VGND sg13g2_fill_1
X_12698_ VGND VPWR _06503_ _06504_ _06507_ _06506_ sg13g2_a21oi_1
X_11718_ _05621_ _05592_ _05620_ _05622_ VPWR VGND sg13g2_nand3_1
XFILLER_30_643 VPWR VGND sg13g2_decap_8
XFILLER_30_654 VPWR VGND sg13g2_decap_8
X_14437_ _00238_ VGND VPWR _00976_ fpmul.seg_reg0.q\[22\] clknet_leaf_93_clk sg13g2_dfrbpq_1
X_11649_ _05498_ _05417_ _05553_ _05554_ VPWR VGND sg13g2_nand3_1
XFILLER_30_676 VPWR VGND sg13g2_fill_2
X_14368_ _00169_ VGND VPWR net1955 fpmul.reg1en.q\[0\] clknet_leaf_95_clk sg13g2_dfrbpq_2
XFILLER_116_737 VPWR VGND sg13g2_decap_8
XFILLER_115_203 VPWR VGND sg13g2_decap_8
X_14299_ _00100_ VGND VPWR _00843_ acc\[9\] clknet_leaf_48_clk sg13g2_dfrbpq_2
XFILLER_124_781 VPWR VGND sg13g2_decap_8
X_08860_ VGND VPWR _03036_ _03038_ _03047_ _03041_ sg13g2_a21oi_1
XFILLER_123_280 VPWR VGND sg13g2_decap_8
XFILLER_112_943 VPWR VGND sg13g2_decap_8
XFILLER_111_420 VPWR VGND sg13g2_fill_1
XFILLER_97_643 VPWR VGND sg13g2_decap_8
X_07811_ _02109_ _02108_ net1640 VPWR VGND sg13g2_nand2_1
XFILLER_97_665 VPWR VGND sg13g2_fill_2
XFILLER_69_345 VPWR VGND sg13g2_decap_8
XFILLER_28_0 VPWR VGND sg13g2_decap_8
X_08791_ _02974_ _02977_ _02978_ VPWR VGND sg13g2_nor2_1
XFILLER_96_164 VPWR VGND sg13g2_decap_4
XFILLER_84_337 VPWR VGND sg13g2_decap_8
X_07742_ _01747_ _02015_ _02047_ VPWR VGND sg13g2_nor2_1
XFILLER_84_359 VPWR VGND sg13g2_decap_8
XFILLER_84_348 VPWR VGND sg13g2_fill_1
XFILLER_38_754 VPWR VGND sg13g2_fill_1
XFILLER_26_905 VPWR VGND sg13g2_decap_8
X_07673_ _01983_ net1793 net1649 acc_sub.exp_mant_logic0.a\[4\] _01949_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_65_562 VPWR VGND sg13g2_decap_8
XFILLER_37_253 VPWR VGND sg13g2_fill_2
XFILLER_80_543 VPWR VGND sg13g2_fill_2
XFILLER_53_746 VPWR VGND sg13g2_fill_1
X_09412_ net1738 _03465_ _03556_ _03557_ VPWR VGND sg13g2_nand3_1
XFILLER_16_28 VPWR VGND sg13g2_decap_8
X_09343_ VGND VPWR _03382_ _03387_ _03495_ _03381_ sg13g2_a21oi_1
XFILLER_61_790 VPWR VGND sg13g2_decap_8
XFILLER_34_982 VPWR VGND sg13g2_decap_8
X_09274_ VPWR _03428_ _03393_ VGND sg13g2_inv_1
XFILLER_20_120 VPWR VGND sg13g2_decap_4
XFILLER_21_643 VPWR VGND sg13g2_fill_2
X_08225_ _02479_ net1645 fp16_sum_pipe.exp_mant_logic0.b\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_32_49 VPWR VGND sg13g2_decap_8
X_08156_ _02414_ _02415_ _02416_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_197 VPWR VGND sg13g2_decap_8
XFILLER_106_203 VPWR VGND sg13g2_fill_1
XFILLER_107_759 VPWR VGND sg13g2_decap_4
XFILLER_106_247 VPWR VGND sg13g2_decap_8
XFILLER_106_7 VPWR VGND sg13g2_decap_8
XFILLER_121_217 VPWR VGND sg13g2_decap_8
XFILLER_115_781 VPWR VGND sg13g2_decap_8
XFILLER_103_932 VPWR VGND sg13g2_decap_8
XFILLER_0_547 VPWR VGND sg13g2_decap_4
XFILLER_114_291 VPWR VGND sg13g2_decap_8
XFILLER_88_687 VPWR VGND sg13g2_decap_8
XFILLER_87_153 VPWR VGND sg13g2_decap_8
XFILLER_48_507 VPWR VGND sg13g2_fill_2
X_08989_ VPWR _03175_ _03173_ VGND sg13g2_inv_1
XFILLER_75_315 VPWR VGND sg13g2_decap_8
XFILLER_87_197 VPWR VGND sg13g2_fill_1
XFILLER_17_905 VPWR VGND sg13g2_decap_8
XFILLER_113_63 VPWR VGND sg13g2_decap_8
XFILLER_90_329 VPWR VGND sg13g2_fill_2
XFILLER_84_860 VPWR VGND sg13g2_fill_2
XFILLER_56_551 VPWR VGND sg13g2_fill_1
XFILLER_44_713 VPWR VGND sg13g2_fill_2
X_10951_ _03586_ _04956_ _04957_ VPWR VGND sg13g2_nor2_1
XFILLER_83_392 VPWR VGND sg13g2_fill_1
X_13670_ VPWR _00221_ net122 VGND sg13g2_inv_1
XFILLER_71_521 VPWR VGND sg13g2_decap_8
XFILLER_56_595 VPWR VGND sg13g2_decap_8
XFILLER_16_426 VPWR VGND sg13g2_fill_1
X_12621_ _06436_ VPWR _06437_ VGND _06421_ fpdiv.div_out\[8\] sg13g2_o21ai_1
XFILLER_73_89 VPWR VGND sg13g2_fill_1
X_10882_ _04893_ _04852_ _04818_ VPWR VGND sg13g2_nand2_1
XFILLER_32_908 VPWR VGND sg13g2_decap_8
XFILLER_43_289 VPWR VGND sg13g2_decap_8
XFILLER_12_621 VPWR VGND sg13g2_decap_8
XFILLER_24_470 VPWR VGND sg13g2_decap_8
XFILLER_106_1013 VPWR VGND sg13g2_fill_1
X_12552_ VGND VPWR _06360_ net1735 _06369_ _06368_ sg13g2_a21oi_1
X_12483_ _06321_ _06185_ _06249_ VPWR VGND sg13g2_nand2_1
XFILLER_40_985 VPWR VGND sg13g2_decap_8
XFILLER_8_614 VPWR VGND sg13g2_decap_8
X_11503_ VGND VPWR _04465_ fp16_sum_pipe.add_renorm0.mantisa\[4\] _05408_ _05407_
+ sg13g2_a21oi_1
X_11434_ _05366_ acc_sub.x2\[10\] net1937 VPWR VGND sg13g2_nand2_1
X_14222_ _00023_ VGND VPWR _00773_ sipo.shift_reg\[3\] clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_7_168 VPWR VGND sg13g2_decap_4
X_14153_ VPWR _00704_ net134 VGND sg13g2_inv_1
XFILLER_98_31 VPWR VGND sg13g2_decap_8
X_11365_ _05317_ _05316_ _05256_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_100_clk clknet_5_15__leaf_clk clknet_leaf_100_clk VPWR VGND sg13g2_buf_8
XFILLER_4_853 VPWR VGND sg13g2_decap_8
X_14084_ VPWR _00635_ net86 VGND sg13g2_inv_1
X_13104_ _06802_ net1700 _06862_ _06863_ VPWR VGND sg13g2_nand3_1
X_11296_ _05255_ _05253_ _05124_ net1697 net1811 VPWR VGND sg13g2_a22oi_1
X_10316_ _04375_ VPWR _01183_ VGND net1919 _04034_ sg13g2_o21ai_1
XFILLER_106_792 VPWR VGND sg13g2_fill_1
XFILLER_79_621 VPWR VGND sg13g2_fill_1
XFILLER_3_385 VPWR VGND sg13g2_decap_8
X_10247_ _04319_ fp16_res_pipe.exp_mant_logic0.b\[1\] net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[4\]
+ _03988_ VPWR VGND sg13g2_a22oi_1
XFILLER_26_1003 VPWR VGND sg13g2_decap_8
XFILLER_79_676 VPWR VGND sg13g2_decap_8
XFILLER_121_784 VPWR VGND sg13g2_decap_8
XFILLER_94_635 VPWR VGND sg13g2_decap_8
XFILLER_79_698 VPWR VGND sg13g2_decap_8
XFILLER_21_7 VPWR VGND sg13g2_decap_8
X_10178_ _03609_ _04222_ _04257_ VPWR VGND sg13g2_nor2_1
XFILLER_94_646 VPWR VGND sg13g2_fill_1
XFILLER_19_220 VPWR VGND sg13g2_decap_4
XFILLER_47_573 VPWR VGND sg13g2_fill_2
X_13937_ VPWR _00488_ net12 VGND sg13g2_inv_1
XFILLER_74_370 VPWR VGND sg13g2_decap_4
XFILLER_35_735 VPWR VGND sg13g2_decap_8
XFILLER_90_885 VPWR VGND sg13g2_fill_1
X_13868_ VPWR _00419_ net50 VGND sg13g2_inv_1
XFILLER_23_919 VPWR VGND sg13g2_decap_8
XFILLER_90_896 VPWR VGND sg13g2_decap_8
X_12819_ _06602_ _06601_ net1732 VPWR VGND sg13g2_nand2_1
X_13799_ VPWR _00350_ net73 VGND sg13g2_inv_1
XFILLER_62_598 VPWR VGND sg13g2_decap_8
XFILLER_31_963 VPWR VGND sg13g2_decap_8
XFILLER_30_451 VPWR VGND sg13g2_fill_2
XFILLER_30_473 VPWR VGND sg13g2_decap_8
XFILLER_8_84 VPWR VGND sg13g2_decap_8
XFILLER_30_484 VPWR VGND sg13g2_fill_2
XFILLER_116_556 VPWR VGND sg13g2_decap_8
XFILLER_104_729 VPWR VGND sg13g2_decap_8
XFILLER_89_418 VPWR VGND sg13g2_decap_8
X_09961_ net1766 net1689 _04056_ VPWR VGND sg13g2_nor2_2
X_08912_ _03009_ _03098_ _03099_ VPWR VGND sg13g2_nor2_2
XFILLER_103_239 VPWR VGND sg13g2_fill_1
XFILLER_100_902 VPWR VGND sg13g2_decap_8
XFILLER_98_974 VPWR VGND sg13g2_decap_8
XFILLER_85_602 VPWR VGND sg13g2_decap_8
X_08843_ VGND VPWR net1788 _03025_ _03030_ _03029_ sg13g2_a21oi_1
XFILLER_111_261 VPWR VGND sg13g2_decap_4
XFILLER_97_473 VPWR VGND sg13g2_fill_2
XFILLER_84_101 VPWR VGND sg13g2_decap_8
XFILLER_57_304 VPWR VGND sg13g2_fill_1
XFILLER_100_979 VPWR VGND sg13g2_decap_8
X_08774_ _02962_ VPWR _01312_ VGND net1899 _02961_ sg13g2_o21ai_1
XFILLER_73_819 VPWR VGND sg13g2_fill_2
X_07725_ _02031_ _01959_ acc_sub.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_38_551 VPWR VGND sg13g2_fill_2
XFILLER_26_702 VPWR VGND sg13g2_decap_8
XFILLER_27_49 VPWR VGND sg13g2_decap_8
XFILLER_25_223 VPWR VGND sg13g2_decap_4
X_07656_ _01967_ net1793 net1646 _01869_ _01935_ VPWR VGND sg13g2_a22oi_1
XFILLER_53_554 VPWR VGND sg13g2_decap_8
XFILLER_25_234 VPWR VGND sg13g2_fill_2
X_07587_ _01832_ net1687 _01901_ VPWR VGND sg13g2_nor2_1
XFILLER_40_226 VPWR VGND sg13g2_fill_2
X_09326_ _03478_ _03477_ _03446_ _03479_ VPWR VGND sg13g2_a21o_1
XFILLER_21_440 VPWR VGND sg13g2_decap_8
X_09257_ VPWR _03411_ _03410_ VGND sg13g2_inv_1
XFILLER_22_996 VPWR VGND sg13g2_decap_8
XFILLER_21_484 VPWR VGND sg13g2_decap_8
XFILLER_21_495 VPWR VGND sg13g2_fill_1
X_08208_ VPWR _02464_ fp16_sum_pipe.exp_mant_logic0.b\[13\] VGND sg13g2_inv_1
X_09188_ _03348_ VPWR _01284_ VGND net1902 _03347_ sg13g2_o21ai_1
XFILLER_4_105 VPWR VGND sg13g2_decap_8
XFILLER_107_545 VPWR VGND sg13g2_fill_1
X_08139_ _02398_ _02399_ _02400_ VPWR VGND sg13g2_nor2b_1
XFILLER_122_515 VPWR VGND sg13g2_fill_2
X_11150_ VPWR _05120_ _05119_ VGND sg13g2_inv_1
XFILLER_108_74 VPWR VGND sg13g2_fill_2
Xplace1880 fpmul.reg1en.q\[0\] net1880 VPWR VGND sg13g2_buf_1
X_10101_ _04182_ _04183_ _04184_ _04185_ VPWR VGND sg13g2_nor3_1
Xplace1891 net1889 net1891 VPWR VGND sg13g2_buf_2
XFILLER_68_67 VPWR VGND sg13g2_decap_8
X_11081_ _05057_ _05049_ acc_sum.exp_mant_logic0.b\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_0_344 VPWR VGND sg13g2_decap_8
XFILLER_1_878 VPWR VGND sg13g2_decap_8
XFILLER_75_101 VPWR VGND sg13g2_decap_8
XFILLER_68_89 VPWR VGND sg13g2_fill_1
XFILLER_48_326 VPWR VGND sg13g2_decap_8
XFILLER_48_304 VPWR VGND sg13g2_fill_2
X_10032_ VPWR _04120_ _04119_ VGND sg13g2_inv_1
XFILLER_76_646 VPWR VGND sg13g2_decap_8
XFILLER_76_657 VPWR VGND sg13g2_fill_2
X_14840_ _00641_ VGND VPWR _01364_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[2\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_1
XFILLER_124_84 VPWR VGND sg13g2_decap_8
X_14771_ _00572_ VGND VPWR _01295_ acc_sub.y\[0\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_29_562 VPWR VGND sg13g2_decap_8
X_13722_ VPWR _00273_ net138 VGND sg13g2_inv_1
XFILLER_91_649 VPWR VGND sg13g2_fill_1
XFILLER_72_841 VPWR VGND sg13g2_fill_2
X_11983_ _05837_ fpmul.reg_a_out\[8\] fpmul.reg_b_out\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_16_201 VPWR VGND sg13g2_fill_2
XFILLER_17_724 VPWR VGND sg13g2_decap_8
XFILLER_17_746 VPWR VGND sg13g2_decap_8
XFILLER_56_1007 VPWR VGND sg13g2_decap_8
X_10934_ VGND VPWR _04845_ _04836_ _04941_ _04739_ sg13g2_a21oi_1
XFILLER_72_896 VPWR VGND sg13g2_fill_2
X_13653_ VPWR _00204_ net70 VGND sg13g2_inv_1
X_10865_ VGND VPWR _04789_ net1825 _04877_ _04876_ sg13g2_a21oi_1
XFILLER_32_727 VPWR VGND sg13g2_decap_8
X_13584_ VPWR _00135_ net118 VGND sg13g2_inv_1
X_12604_ _06399_ _06401_ _06420_ VPWR VGND sg13g2_xor2_1
X_12535_ _06353_ VPWR _00942_ VGND net1957 _05891_ sg13g2_o21ai_1
XFILLER_40_771 VPWR VGND sg13g2_fill_2
XFILLER_8_411 VPWR VGND sg13g2_decap_8
XFILLER_9_934 VPWR VGND sg13g2_decap_8
XFILLER_13_996 VPWR VGND sg13g2_decap_8
X_10796_ VGND VPWR _04807_ _04808_ _04806_ _04775_ sg13g2_a21oi_2
XFILLER_33_70 VPWR VGND sg13g2_decap_8
XFILLER_33_92 VPWR VGND sg13g2_decap_8
XFILLER_69_7 VPWR VGND sg13g2_decap_8
X_12466_ _06308_ _06307_ _06305_ VPWR VGND sg13g2_nand2b_1
X_14205_ VPWR _00756_ net99 VGND sg13g2_inv_1
X_11417_ _05355_ net1647 net1718 VPWR VGND sg13g2_nand2_1
X_12397_ _06243_ _06187_ _06188_ VPWR VGND sg13g2_nand2_1
XFILLER_126_876 VPWR VGND sg13g2_decap_8
XFILLER_125_342 VPWR VGND sg13g2_fill_1
XFILLER_113_515 VPWR VGND sg13g2_fill_1
XFILLER_98_204 VPWR VGND sg13g2_decap_8
X_14136_ VPWR _00687_ net114 VGND sg13g2_inv_1
X_11348_ _05301_ _05211_ _05253_ VPWR VGND sg13g2_nand2_1
X_14067_ VPWR _00618_ net95 VGND sg13g2_inv_1
X_11279_ _05241_ net1761 acc_sum.op_sign_logic0.mantisa_a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_3_182 VPWR VGND sg13g2_decap_8
X_13018_ _06785_ VPWR _06786_ VGND net1853 fpmul.seg_reg0.q\[10\] sg13g2_o21ai_1
XFILLER_79_462 VPWR VGND sg13g2_fill_2
XFILLER_79_495 VPWR VGND sg13g2_decap_8
XFILLER_39_348 VPWR VGND sg13g2_fill_1
XFILLER_95_988 VPWR VGND sg13g2_decap_8
XFILLER_55_819 VPWR VGND sg13g2_decap_8
X_14969_ _00770_ VGND VPWR _01489_ acc_sub.seg_reg1.q\[21\] clknet_leaf_42_clk sg13g2_dfrbpq_2
X_07510_ VPWR _01832_ _01831_ VGND sg13g2_inv_1
XFILLER_35_532 VPWR VGND sg13g2_decap_8
X_08490_ _02718_ fpdiv.divider0.remainder_reg\[6\] net1708 net1748 fpdiv.divider0.dividend\[6\]
+ VPWR VGND sg13g2_a22oi_1
X_07441_ _01771_ net1749 fpdiv.divider0.divisor\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_63_896 VPWR VGND sg13g2_fill_1
Xfanout19 net24 net19 VPWR VGND sg13g2_buf_2
XFILLER_50_513 VPWR VGND sg13g2_decap_8
XFILLER_35_587 VPWR VGND sg13g2_decap_4
XFILLER_95_0 VPWR VGND sg13g2_decap_8
X_07372_ _01723_ acc\[15\] VPWR VGND sg13g2_inv_2
XFILLER_16_790 VPWR VGND sg13g2_decap_8
X_09111_ _03135_ _03292_ _03290_ _03293_ VPWR VGND sg13g2_nand3_1
XFILLER_31_760 VPWR VGND sg13g2_fill_1
X_09042_ _03228_ _03227_ acc_sub.add_renorm0.exp\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_117_865 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
X_09944_ _04040_ _04039_ _04009_ VPWR VGND sg13g2_nand2_1
XFILLER_112_570 VPWR VGND sg13g2_decap_8
X_09875_ VGND VPWR _03979_ net1820 _01229_ _03980_ sg13g2_a21oi_1
XFILLER_98_782 VPWR VGND sg13g2_decap_8
X_08826_ _03013_ _02990_ VPWR VGND sg13g2_inv_2
XFILLER_112_581 VPWR VGND sg13g2_fill_2
XFILLER_86_966 VPWR VGND sg13g2_decap_8
XFILLER_57_134 VPWR VGND sg13g2_decap_8
XFILLER_46_808 VPWR VGND sg13g2_decap_8
X_08757_ _02951_ acc_sum.exp_mant_logic0.a\[6\] VPWR VGND sg13g2_inv_2
XFILLER_73_649 VPWR VGND sg13g2_decap_4
XFILLER_57_189 VPWR VGND sg13g2_decap_8
XFILLER_54_14 VPWR VGND sg13g2_decap_8
XFILLER_39_882 VPWR VGND sg13g2_decap_8
X_07708_ _02015_ _01989_ VPWR VGND sg13g2_inv_2
X_08688_ VGND VPWR net1671 _02847_ _02903_ net1739 sg13g2_a21oi_1
XFILLER_72_159 VPWR VGND sg13g2_fill_2
X_07639_ _01952_ net1646 _01869_ VPWR VGND sg13g2_nand2_1
XFILLER_14_738 VPWR VGND sg13g2_fill_1
XFILLER_110_42 VPWR VGND sg13g2_decap_8
XFILLER_13_226 VPWR VGND sg13g2_fill_2
XFILLER_14_749 VPWR VGND sg13g2_fill_1
X_09309_ _03462_ _03461_ _03407_ VPWR VGND sg13g2_nand2b_1
XFILLER_9_219 VPWR VGND sg13g2_fill_2
X_10581_ _04603_ VPWR _01146_ VGND net1930 _02208_ sg13g2_o21ai_1
XFILLER_10_933 VPWR VGND sg13g2_decap_8
XFILLER_127_629 VPWR VGND sg13g2_decap_8
XFILLER_127_618 VPWR VGND sg13g2_decap_8
XFILLER_108_810 VPWR VGND sg13g2_fill_2
X_12320_ _06065_ _06165_ _06166_ VPWR VGND sg13g2_nor2_1
X_12251_ _05962_ _05961_ _05956_ _06097_ VPWR VGND sg13g2_nand3_1
XFILLER_6_948 VPWR VGND sg13g2_decap_8
XFILLER_5_436 VPWR VGND sg13g2_decap_8
XFILLER_123_813 VPWR VGND sg13g2_decap_8
XFILLER_119_84 VPWR VGND sg13g2_decap_8
X_11202_ _05169_ _05075_ acc_sum.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
X_12182_ VPWR _06028_ _06027_ VGND sg13g2_inv_1
XFILLER_89_760 VPWR VGND sg13g2_decap_8
X_11133_ VGND VPWR _05090_ _05048_ _05103_ _05102_ sg13g2_a21oi_1
XFILLER_1_653 VPWR VGND sg13g2_decap_8
XFILLER_95_32 VPWR VGND sg13g2_decap_8
XFILLER_77_911 VPWR VGND sg13g2_fill_1
X_11064_ _05042_ _05035_ _05041_ VPWR VGND sg13g2_nand2_2
XFILLER_49_624 VPWR VGND sg13g2_fill_2
XFILLER_95_43 VPWR VGND sg13g2_fill_1
XFILLER_77_955 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
X_10015_ _04100_ _04102_ _04103_ VPWR VGND sg13g2_nor2_1
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_91_446 VPWR VGND sg13g2_decap_8
XFILLER_91_435 VPWR VGND sg13g2_decap_8
X_14823_ _00624_ VGND VPWR _01347_ acc_sum.seg_reg1.q\[20\] clknet_leaf_24_clk sg13g2_dfrbpq_1
XFILLER_76_487 VPWR VGND sg13g2_decap_8
XFILLER_63_104 VPWR VGND sg13g2_fill_1
XFILLER_48_189 VPWR VGND sg13g2_fill_1
XFILLER_28_70 VPWR VGND sg13g2_decap_8
XFILLER_91_457 VPWR VGND sg13g2_decap_8
X_14754_ _00555_ VGND VPWR net1899 acc_sum.reg1en.q\[0\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_11966_ VPWR _05821_ fpmul.seg_reg0.q\[24\] VGND sg13g2_inv_1
XFILLER_17_532 VPWR VGND sg13g2_fill_2
XFILLER_17_543 VPWR VGND sg13g2_fill_1
X_13705_ VPWR _00256_ net65 VGND sg13g2_inv_1
XFILLER_45_896 VPWR VGND sg13g2_decap_4
X_10917_ net1771 VPWR _04926_ VGND _04875_ _04925_ sg13g2_o21ai_1
X_14685_ _00486_ VGND VPWR _01213_ fp16_res_pipe.seg_reg0.q\[22\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_1
XFILLER_71_192 VPWR VGND sg13g2_decap_8
X_13636_ VPWR _00187_ net85 VGND sg13g2_inv_1
X_11897_ fpmul.seg_reg0.q\[51\] fpmul.reg_a_out\[12\] net1878 _01005_ VPWR VGND sg13g2_mux2_1
XFILLER_44_91 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_fill_1
X_10848_ VGND VPWR _04814_ net1825 _04860_ _04859_ sg13g2_a21oi_1
XFILLER_81_6 VPWR VGND sg13g2_fill_1
X_13567_ VPWR _00118_ net33 VGND sg13g2_inv_1
XFILLER_8_230 VPWR VGND sg13g2_decap_4
X_10779_ _04790_ VPWR _04791_ VGND _04786_ _04789_ sg13g2_o21ai_1
X_13498_ VPWR _00049_ net33 VGND sg13g2_inv_1
X_12518_ VGND VPWR _03601_ net1955 _00950_ _06344_ sg13g2_a21oi_1
XFILLER_9_764 VPWR VGND sg13g2_decap_8
X_12449_ _06288_ _06283_ _06294_ VPWR VGND sg13g2_nor2_1
XFILLER_8_274 VPWR VGND sg13g2_fill_2
XFILLER_125_161 VPWR VGND sg13g2_decap_8
XFILLER_114_846 VPWR VGND sg13g2_decap_8
XFILLER_113_312 VPWR VGND sg13g2_fill_2
XFILLER_5_63 VPWR VGND sg13g2_decap_8
XFILLER_99_557 VPWR VGND sg13g2_fill_1
X_07990_ _02258_ fp16_sum_pipe.exp_mant_logic0.a\[7\] _02250_ fp16_sum_pipe.seg_reg0.q\[22\]
+ net1775 VPWR VGND sg13g2_a22oi_1
X_14119_ VPWR _00670_ net43 VGND sg13g2_inv_1
X_09660_ _03777_ _03674_ _03666_ _03655_ _03630_ VPWR VGND sg13g2_a22oi_1
XFILLER_95_752 VPWR VGND sg13g2_fill_2
XFILLER_95_730 VPWR VGND sg13g2_decap_4
XFILLER_79_292 VPWR VGND sg13g2_decap_8
XFILLER_79_281 VPWR VGND sg13g2_fill_1
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_94_240 VPWR VGND sg13g2_decap_8
XFILLER_94_251 VPWR VGND sg13g2_fill_2
X_08611_ _02833_ VPWR _02834_ VGND _02813_ _02832_ sg13g2_o21ai_1
XFILLER_83_925 VPWR VGND sg13g2_decap_8
XFILLER_55_605 VPWR VGND sg13g2_decap_8
XFILLER_10_0 VPWR VGND sg13g2_decap_8
X_09591_ net1805 acc_sum.add_renorm0.mantisa\[2\] _03708_ VPWR VGND sg13g2_nor2_1
XFILLER_27_318 VPWR VGND sg13g2_decap_8
X_08542_ VGND VPWR _02760_ _02762_ _02766_ _02765_ sg13g2_a21oi_1
XFILLER_70_619 VPWR VGND sg13g2_decap_8
XFILLER_36_863 VPWR VGND sg13g2_fill_1
XFILLER_35_340 VPWR VGND sg13g2_fill_1
X_08473_ _02703_ VPWR _02704_ VGND fpdiv.divider0.remainder_reg\[8\] net1647 sg13g2_o21ai_1
XFILLER_36_885 VPWR VGND sg13g2_decap_8
XFILLER_35_373 VPWR VGND sg13g2_decap_8
X_07424_ VPWR _01759_ fpdiv.divider0.divisor_reg\[11\] VGND sg13g2_inv_1
XFILLER_90_490 VPWR VGND sg13g2_decap_8
XFILLER_62_192 VPWR VGND sg13g2_decap_8
XFILLER_24_28 VPWR VGND sg13g2_decap_8
XFILLER_11_719 VPWR VGND sg13g2_decap_8
X_07355_ _01712_ VPWR _01474_ VGND net1797 _01711_ sg13g2_o21ai_1
XFILLER_10_229 VPWR VGND sg13g2_decap_8
X_07286_ _01653_ VPWR _01654_ VGND _01507_ _01652_ sg13g2_o21ai_1
X_09025_ _03211_ _03210_ _03198_ VPWR VGND sg13g2_nand2_1
XFILLER_108_139 VPWR VGND sg13g2_decap_8
XFILLER_40_49 VPWR VGND sg13g2_decap_8
XFILLER_117_662 VPWR VGND sg13g2_fill_1
XFILLER_104_301 VPWR VGND sg13g2_decap_8
XFILLER_116_194 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_120_827 VPWR VGND sg13g2_decap_8
XFILLER_104_389 VPWR VGND sg13g2_fill_2
X_09927_ _04024_ _03599_ fp16_res_pipe.exp_mant_logic0.b\[9\] VPWR VGND sg13g2_nand2_2
XFILLER_105_75 VPWR VGND sg13g2_decap_4
X_09858_ _03733_ _03807_ _03967_ VPWR VGND sg13g2_xor2_1
XFILLER_100_540 VPWR VGND sg13g2_decap_4
XFILLER_59_999 VPWR VGND sg13g2_fill_1
X_08809_ _02996_ _02982_ _02976_ VPWR VGND sg13g2_xnor2_1
XFILLER_100_595 VPWR VGND sg13g2_decap_8
X_09789_ _03903_ _03818_ _03799_ VPWR VGND sg13g2_nand2_1
XFILLER_74_947 VPWR VGND sg13g2_fill_1
XFILLER_65_35 VPWR VGND sg13g2_decap_8
XFILLER_58_487 VPWR VGND sg13g2_fill_1
XFILLER_46_638 VPWR VGND sg13g2_fill_2
XFILLER_45_126 VPWR VGND sg13g2_decap_8
XFILLER_74_969 VPWR VGND sg13g2_fill_1
XFILLER_73_446 VPWR VGND sg13g2_fill_2
X_11820_ VGND VPWR _05720_ _05638_ _05639_ sg13g2_or2_1
XFILLER_73_479 VPWR VGND sg13g2_fill_2
X_11751_ net1839 _04587_ _05655_ VPWR VGND sg13g2_nor2_1
XFILLER_121_63 VPWR VGND sg13g2_decap_8
XFILLER_81_23 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_80_clk clknet_5_26__leaf_clk clknet_leaf_80_clk VPWR VGND sg13g2_buf_8
XFILLER_53_170 VPWR VGND sg13g2_decap_8
XFILLER_41_332 VPWR VGND sg13g2_fill_1
X_10702_ VPWR _04715_ _04714_ VGND sg13g2_inv_1
X_14470_ _00271_ VGND VPWR _01009_ fpdiv.divider0.counter\[0\] clknet_leaf_71_clk
+ sg13g2_dfrbpq_1
X_11682_ _04581_ net1727 _05586_ VPWR VGND sg13g2_nor2_1
X_13421_ _07089_ VPWR _00793_ VGND _07046_ net1720 sg13g2_o21ai_1
X_10633_ _04613_ _04645_ _04646_ VPWR VGND sg13g2_nor2_1
X_13352_ _07050_ net1723 fp16_res_pipe.x2\[4\] VPWR VGND sg13g2_nand2_1
X_10564_ _04594_ VPWR _01154_ VGND net1844 _04593_ sg13g2_o21ai_1
XFILLER_127_426 VPWR VGND sg13g2_decap_8
X_12303_ _06141_ _06143_ _06149_ VPWR VGND sg13g2_xor2_1
XFILLER_6_723 VPWR VGND sg13g2_fill_2
X_13283_ _06999_ sipo.word\[6\] VPWR VGND sg13g2_inv_2
X_10495_ _04384_ VPWR _04540_ VGND _04539_ net1673 sg13g2_o21ai_1
X_12234_ _06080_ net1859 net1866 VPWR VGND sg13g2_nand2_1
X_12165_ _06009_ _06010_ _05981_ _06011_ VPWR VGND sg13g2_nand3_1
XFILLER_2_940 VPWR VGND sg13g2_decap_8
XFILLER_122_175 VPWR VGND sg13g2_decap_8
XFILLER_111_838 VPWR VGND sg13g2_decap_8
XFILLER_96_527 VPWR VGND sg13g2_decap_8
X_11116_ VGND VPWR _05085_ _05038_ _05086_ _05000_ sg13g2_a21oi_1
XFILLER_7_1000 VPWR VGND sg13g2_decap_8
XFILLER_1_450 VPWR VGND sg13g2_decap_8
XFILLER_77_741 VPWR VGND sg13g2_fill_1
X_12096_ _05888_ _05886_ _05941_ _05942_ VPWR VGND sg13g2_nand3_1
XFILLER_49_432 VPWR VGND sg13g2_fill_1
XFILLER_49_410 VPWR VGND sg13g2_fill_2
X_11047_ _05026_ _05011_ _05025_ VPWR VGND sg13g2_nand2_2
XFILLER_65_914 VPWR VGND sg13g2_decap_8
XFILLER_49_443 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_92_733 VPWR VGND sg13g2_decap_8
XFILLER_76_295 VPWR VGND sg13g2_decap_4
X_14806_ _00607_ VGND VPWR _01330_ acc_sum.add_renorm0.exp\[3\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
XFILLER_91_232 VPWR VGND sg13g2_decap_8
XFILLER_64_468 VPWR VGND sg13g2_decap_8
XFILLER_92_788 VPWR VGND sg13g2_fill_1
X_12998_ fpmul.seg_reg0.q\[15\] fpmul.seg_reg0.q\[14\] _06766_ VPWR VGND sg13g2_nor2_1
XFILLER_45_671 VPWR VGND sg13g2_decap_8
XFILLER_18_885 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_71_clk clknet_5_31__leaf_clk clknet_leaf_71_clk VPWR VGND sg13g2_buf_8
X_11949_ _05810_ net1884 net1863 VPWR VGND sg13g2_nand2_1
XFILLER_44_192 VPWR VGND sg13g2_fill_1
X_14737_ _00538_ VGND VPWR _01265_ fp16_res_pipe.add_renorm0.mantisa\[0\] clknet_leaf_137_clk
+ sg13g2_dfrbpq_1
X_14668_ _00469_ VGND VPWR _01196_ fp16_res_pipe.op_sign_logic0.mantisa_b\[5\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_2
XFILLER_119_905 VPWR VGND sg13g2_decap_8
X_13619_ VPWR _00170_ net65 VGND sg13g2_inv_1
XFILLER_20_549 VPWR VGND sg13g2_fill_1
XFILLER_118_404 VPWR VGND sg13g2_decap_8
X_07140_ VPWR _01512_ _01511_ VGND sg13g2_inv_1
XFILLER_72_2 VPWR VGND sg13g2_fill_1
X_14599_ _00400_ VGND VPWR _01131_ fp16_res_pipe.y\[10\] clknet_leaf_129_clk sg13g2_dfrbpq_1
XFILLER_9_583 VPWR VGND sg13g2_fill_2
XFILLER_127_960 VPWR VGND sg13g2_decap_8
XFILLER_58_0 VPWR VGND sg13g2_decap_8
XFILLER_114_654 VPWR VGND sg13g2_fill_2
XFILLER_114_643 VPWR VGND sg13g2_decap_8
XFILLER_102_827 VPWR VGND sg13g2_fill_1
X_09712_ _03642_ acc_sum.add_renorm0.mantisa\[10\] _03828_ VPWR VGND sg13g2_nor2b_2
XFILLER_68_730 VPWR VGND sg13g2_decap_8
XFILLER_19_28 VPWR VGND sg13g2_decap_8
X_07973_ _02179_ _02245_ _02246_ VPWR VGND sg13g2_nor2_2
XFILLER_110_871 VPWR VGND sg13g2_decap_8
XFILLER_101_359 VPWR VGND sg13g2_decap_8
XFILLER_68_763 VPWR VGND sg13g2_decap_4
X_09643_ _03760_ _03649_ _03674_ VPWR VGND sg13g2_nand2_1
XFILLER_95_593 VPWR VGND sg13g2_decap_8
XFILLER_67_273 VPWR VGND sg13g2_decap_8
X_09574_ _03690_ VPWR _03691_ VGND net1806 _03620_ sg13g2_o21ai_1
XFILLER_55_468 VPWR VGND sg13g2_decap_8
X_08525_ VPWR _02749_ acc_sum.op_sign_logic0.mantisa_a\[3\] VGND sg13g2_inv_1
XFILLER_35_49 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_62_clk clknet_5_28__leaf_clk clknet_leaf_62_clk VPWR VGND sg13g2_buf_8
X_08456_ VPWR _02689_ fpdiv.divider0.remainder_reg\[11\] VGND sg13g2_inv_1
XFILLER_50_140 VPWR VGND sg13g2_decap_8
XFILLER_23_354 VPWR VGND sg13g2_decap_8
X_07407_ _01746_ VPWR _01456_ VGND net1889 _01745_ sg13g2_o21ai_1
X_08387_ _02621_ _02622_ _02620_ _02625_ VPWR VGND _02624_ sg13g2_nand4_1
XFILLER_11_516 VPWR VGND sg13g2_decap_8
X_07338_ _01699_ VPWR _01478_ VGND _01695_ _01696_ sg13g2_o21ai_1
XFILLER_118_971 VPWR VGND sg13g2_decap_8
X_07269_ _01638_ _01513_ _01613_ VPWR VGND sg13g2_nand2b_1
XFILLER_124_429 VPWR VGND sg13g2_fill_1
X_09008_ _03009_ _03157_ _03173_ _03194_ VPWR VGND sg13g2_nor3_1
XFILLER_117_481 VPWR VGND sg13g2_decap_8
X_10280_ _04349_ _04190_ fp16_res_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_104_197 VPWR VGND sg13g2_decap_8
XFILLER_104_186 VPWR VGND sg13g2_fill_1
XFILLER_59_741 VPWR VGND sg13g2_decap_8
XFILLER_59_730 VPWR VGND sg13g2_decap_4
XFILLER_116_96 VPWR VGND sg13g2_decap_8
XFILLER_93_508 VPWR VGND sg13g2_decap_8
X_13970_ VPWR _00521_ net25 VGND sg13g2_inv_1
XFILLER_19_605 VPWR VGND sg13g2_fill_1
X_12921_ acc\[4\] net1907 _03983_ _06695_ VPWR VGND sg13g2_nand3_1
XFILLER_18_115 VPWR VGND sg13g2_decap_4
XFILLER_100_392 VPWR VGND sg13g2_decap_4
XFILLER_74_755 VPWR VGND sg13g2_fill_1
XFILLER_62_917 VPWR VGND sg13g2_fill_2
XFILLER_73_276 VPWR VGND sg13g2_fill_1
X_12852_ _06632_ _06628_ _06631_ _06627_ net1943 VPWR VGND sg13g2_a22oi_1
XFILLER_55_980 VPWR VGND sg13g2_fill_2
XFILLER_92_88 VPWR VGND sg13g2_fill_1
X_12783_ VPWR _06568_ piso.tx_bit_counter\[2\] VGND sg13g2_inv_1
Xclkbuf_leaf_53_clk clknet_5_18__leaf_clk clknet_leaf_53_clk VPWR VGND sg13g2_buf_8
X_11803_ _05656_ VPWR _05704_ VGND _05659_ _05668_ sg13g2_o21ai_1
XFILLER_15_833 VPWR VGND sg13g2_fill_2
X_14522_ _00323_ VGND VPWR _01058_ fpdiv.reg_a_out\[13\] clknet_leaf_126_clk sg13g2_dfrbpq_2
XFILLER_14_365 VPWR VGND sg13g2_decap_8
X_11734_ VGND VPWR _05635_ _05636_ _05638_ _05637_ sg13g2_a21oi_1
X_14453_ _00254_ VGND VPWR _00992_ fpmul.seg_reg0.q\[38\] clknet_leaf_122_clk sg13g2_dfrbpq_1
XFILLER_14_387 VPWR VGND sg13g2_decap_8
X_11665_ _05541_ _05551_ _05516_ _05570_ VPWR VGND _05569_ sg13g2_nand4_1
X_13404_ _07080_ VPWR _00801_ VGND _07026_ net1721 sg13g2_o21ai_1
Xclkbuf_4_6_0_clk clknet_0_clk clknet_4_6_0_clk VPWR VGND sg13g2_buf_8
X_10616_ net1823 fp16_res_pipe.add_renorm0.mantisa\[2\] _04629_ VPWR VGND sg13g2_nor2_1
X_14384_ _00185_ VGND VPWR _00925_ fpmul.reg_b_out\[15\] clknet_leaf_126_clk sg13g2_dfrbpq_1
XFILLER_10_571 VPWR VGND sg13g2_fill_1
X_11596_ _05501_ net1841 fp16_sum_pipe.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_127_245 VPWR VGND sg13g2_decap_8
XFILLER_116_919 VPWR VGND sg13g2_decap_8
X_13335_ _07039_ VPWR _00829_ VGND _07037_ net1726 sg13g2_o21ai_1
XFILLER_41_70 VPWR VGND sg13g2_decap_8
X_10547_ VPWR _04583_ fp16_sum_pipe.add_renorm0.exp\[6\] VGND sg13g2_inv_1
Xplace1709 _04775_ net1709 VPWR VGND sg13g2_buf_2
X_13266_ _03283_ _02576_ _06986_ VPWR VGND sg13g2_nor2_1
XFILLER_51_7 VPWR VGND sg13g2_decap_8
XFILLER_6_586 VPWR VGND sg13g2_fill_1
XFILLER_6_564 VPWR VGND sg13g2_decap_8
X_10478_ _04460_ _04524_ _04525_ VPWR VGND sg13g2_nor2_1
XFILLER_124_963 VPWR VGND sg13g2_decap_8
X_12217_ _06063_ net1856 net1868 VPWR VGND sg13g2_nand2_1
XFILLER_111_613 VPWR VGND sg13g2_fill_2
XFILLER_69_527 VPWR VGND sg13g2_decap_8
X_13197_ _06932_ VPWR _00860_ VGND _06931_ net1713 sg13g2_o21ai_1
XFILLER_123_495 VPWR VGND sg13g2_fill_1
XFILLER_111_635 VPWR VGND sg13g2_decap_8
X_12148_ _05994_ _05992_ _05993_ VPWR VGND sg13g2_nand2_1
X_12079_ _05925_ fpmul.reg_a_out\[6\] net1866 VPWR VGND sg13g2_nand2_1
XFILLER_2_42 VPWR VGND sg13g2_decap_8
XFILLER_110_167 VPWR VGND sg13g2_decap_8
XFILLER_65_733 VPWR VGND sg13g2_fill_2
XFILLER_65_722 VPWR VGND sg13g2_decap_8
XFILLER_38_925 VPWR VGND sg13g2_decap_8
XFILLER_37_457 VPWR VGND sg13g2_decap_4
XFILLER_65_777 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_44_clk clknet_5_23__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
XFILLER_80_747 VPWR VGND sg13g2_fill_2
XFILLER_64_287 VPWR VGND sg13g2_fill_1
XFILLER_18_693 VPWR VGND sg13g2_decap_8
XFILLER_33_663 VPWR VGND sg13g2_fill_2
X_08310_ _02554_ _02555_ _02556_ VPWR VGND _02553_ sg13g2_nand3b_1
X_09290_ VPWR _03444_ fp16_res_pipe.op_sign_logic0.mantisa_a\[10\] VGND sg13g2_inv_1
XFILLER_33_696 VPWR VGND sg13g2_fill_1
X_08241_ _02493_ net1842 _02338_ _02275_ fp16_sum_pipe.exp_mant_logic0.b\[3\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_21_825 VPWR VGND sg13g2_decap_8
XFILLER_20_357 VPWR VGND sg13g2_decap_8
X_08172_ _02425_ _02430_ _02424_ _02431_ VPWR VGND sg13g2_nand3_1
XFILLER_119_779 VPWR VGND sg13g2_decap_8
XFILLER_118_245 VPWR VGND sg13g2_decap_8
X_07123_ net1783 _01495_ _01496_ VPWR VGND sg13g2_nor2_1
XFILLER_9_380 VPWR VGND sg13g2_decap_8
XFILLER_106_407 VPWR VGND sg13g2_fill_2
XFILLER_115_963 VPWR VGND sg13g2_decap_8
XFILLER_82_1003 VPWR VGND sg13g2_decap_8
XFILLER_114_462 VPWR VGND sg13g2_decap_4
XFILLER_88_803 VPWR VGND sg13g2_fill_1
XFILLER_88_869 VPWR VGND sg13g2_decap_4
X_07956_ VPWR _02230_ _02211_ VGND sg13g2_inv_1
XFILLER_96_880 VPWR VGND sg13g2_decap_8
XFILLER_68_582 VPWR VGND sg13g2_decap_4
XFILLER_56_733 VPWR VGND sg13g2_decap_4
XFILLER_95_390 VPWR VGND sg13g2_decap_8
X_07887_ _02170_ VPWR _01400_ VGND net1892 _02096_ sg13g2_o21ai_1
XFILLER_83_530 VPWR VGND sg13g2_decap_4
XFILLER_56_766 VPWR VGND sg13g2_fill_1
XFILLER_56_755 VPWR VGND sg13g2_decap_8
XFILLER_29_969 VPWR VGND sg13g2_decap_8
X_09626_ net1802 _03742_ _03743_ VPWR VGND sg13g2_nor2_1
XFILLER_102_21 VPWR VGND sg13g2_decap_8
XFILLER_56_777 VPWR VGND sg13g2_decap_8
XFILLER_43_405 VPWR VGND sg13g2_fill_2
XFILLER_37_980 VPWR VGND sg13g2_decap_8
XFILLER_15_107 VPWR VGND sg13g2_fill_1
XFILLER_16_619 VPWR VGND sg13g2_fill_1
X_09557_ VGND VPWR _03622_ _03674_ _03673_ _03672_ sg13g2_a21oi_2
XFILLER_71_747 VPWR VGND sg13g2_decap_8
XFILLER_71_736 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_35_clk clknet_5_20__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
X_08508_ _02730_ _02731_ _02732_ VPWR VGND sg13g2_nor2_1
XFILLER_12_803 VPWR VGND sg13g2_decap_8
XFILLER_24_652 VPWR VGND sg13g2_fill_2
X_09488_ _03610_ acc_sub.x2\[4\] net1918 VPWR VGND sg13g2_nand2_1
X_08439_ _02673_ _02671_ _02672_ VPWR VGND sg13g2_nand2_1
XFILLER_11_313 VPWR VGND sg13g2_decap_8
XFILLER_8_807 VPWR VGND sg13g2_fill_2
XFILLER_12_869 VPWR VGND sg13g2_decap_8
X_11450_ VPWR _05376_ fpdiv.divider0.dividend\[8\] VGND sg13g2_inv_1
XFILLER_7_328 VPWR VGND sg13g2_fill_2
X_11381_ _05331_ net1812 _05227_ acc_sum.exp_mant_logic0.b\[4\] _05211_ VPWR VGND
+ sg13g2_a22oi_1
X_10401_ VPWR _04451_ _04397_ VGND sg13g2_inv_1
X_13120_ _06868_ _06779_ _06875_ VPWR VGND sg13g2_xor2_1
X_10332_ _04383_ VPWR _01175_ VGND net1921 _04322_ sg13g2_o21ai_1
X_13051_ _06819_ _06818_ fpmul.seg_reg0.q\[22\] VPWR VGND sg13g2_nand2_1
XFILLER_11_84 VPWR VGND sg13g2_decap_8
XFILLER_127_84 VPWR VGND sg13g2_decap_8
XFILLER_124_259 VPWR VGND sg13g2_decap_8
XFILLER_106_985 VPWR VGND sg13g2_decap_8
X_12002_ _05856_ _05854_ _05855_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_567 VPWR VGND sg13g2_decap_8
X_10263_ _04334_ _04333_ _04272_ VPWR VGND sg13g2_nand2_1
X_10194_ _04271_ net1745 net1644 net1688 net1829 VPWR VGND sg13g2_a22oi_1
XFILLER_121_966 VPWR VGND sg13g2_decap_8
X_13953_ VPWR _00504_ net97 VGND sg13g2_inv_1
XFILLER_47_744 VPWR VGND sg13g2_decap_8
XFILLER_46_232 VPWR VGND sg13g2_decap_8
XFILLER_19_435 VPWR VGND sg13g2_fill_1
XFILLER_19_446 VPWR VGND sg13g2_decap_8
X_12904_ _06680_ _06679_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_59_1005 VPWR VGND sg13g2_decap_8
XFILLER_35_939 VPWR VGND sg13g2_decap_8
X_13884_ VPWR _00435_ net48 VGND sg13g2_inv_1
XFILLER_28_980 VPWR VGND sg13g2_decap_8
X_12835_ VGND VPWR net1935 add_result\[11\] _06616_ net1943 sg13g2_a21oi_1
XFILLER_62_736 VPWR VGND sg13g2_decap_8
XFILLER_61_224 VPWR VGND sg13g2_decap_8
XFILLER_36_70 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_5_16__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_50_909 VPWR VGND sg13g2_fill_1
XFILLER_99_7 VPWR VGND sg13g2_fill_2
XFILLER_70_780 VPWR VGND sg13g2_decap_4
X_14505_ _00306_ VGND VPWR _01041_ fpdiv.reg_b_out\[12\] clknet_leaf_53_clk sg13g2_dfrbpq_2
X_12766_ _06550_ VPWR _06551_ VGND _06546_ div_result\[15\] sg13g2_o21ai_1
XFILLER_15_674 VPWR VGND sg13g2_decap_8
X_12697_ _06454_ _06456_ _06449_ _06506_ VPWR VGND _06505_ sg13g2_nand4_1
XFILLER_42_493 VPWR VGND sg13g2_decap_4
X_11717_ _05621_ _05604_ VPWR VGND sg13g2_inv_2
X_14436_ _00237_ VGND VPWR _00975_ fpmul.seg_reg0.q\[21\] clknet_leaf_96_clk sg13g2_dfrbpq_1
X_11648_ _05553_ _05522_ _05408_ VPWR VGND sg13g2_nand2_1
XFILLER_116_705 VPWR VGND sg13g2_fill_1
X_14367_ _00168_ VGND VPWR _00909_ _00020_ clknet_leaf_86_clk sg13g2_dfrbpq_1
X_11579_ _05477_ _05428_ _05484_ VPWR VGND sg13g2_nor2_1
X_13318_ _07027_ _02563_ sipo.word_ready VPWR VGND sg13g2_nand2_2
XFILLER_7_895 VPWR VGND sg13g2_decap_8
X_14298_ _00099_ VGND VPWR _00842_ acc\[8\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_66_1009 VPWR VGND sg13g2_decap_4
XFILLER_124_760 VPWR VGND sg13g2_decap_8
XFILLER_115_259 VPWR VGND sg13g2_decap_8
XFILLER_97_611 VPWR VGND sg13g2_fill_2
X_13249_ _06973_ net1729 acc_sum.y\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_112_922 VPWR VGND sg13g2_decap_8
XFILLER_69_324 VPWR VGND sg13g2_decap_8
X_08790_ acc_sub.add_renorm0.mantisa\[8\] acc_sub.add_renorm0.mantisa\[7\] _02976_
+ _02977_ VPWR VGND sg13g2_nand3_1
XFILLER_111_443 VPWR VGND sg13g2_decap_4
X_07810_ _02106_ _02107_ _02105_ _02108_ VPWR VGND sg13g2_nand3_1
XFILLER_96_143 VPWR VGND sg13g2_decap_8
XFILLER_112_999 VPWR VGND sg13g2_decap_8
X_07741_ VGND VPWR acc_sub.exp_mant_logic0.a\[2\] _01975_ _02046_ _02045_ sg13g2_a21oi_1
XFILLER_84_316 VPWR VGND sg13g2_decap_8
XFILLER_78_880 VPWR VGND sg13g2_decap_8
XFILLER_69_379 VPWR VGND sg13g2_decap_8
XFILLER_38_711 VPWR VGND sg13g2_decap_8
XFILLER_65_541 VPWR VGND sg13g2_decap_8
XFILLER_37_232 VPWR VGND sg13g2_decap_8
X_07672_ _01982_ _01935_ net1792 VPWR VGND sg13g2_nand2_1
XFILLER_92_360 VPWR VGND sg13g2_fill_1
XFILLER_38_788 VPWR VGND sg13g2_fill_1
XFILLER_38_777 VPWR VGND sg13g2_decap_8
XFILLER_65_585 VPWR VGND sg13g2_decap_8
X_09411_ _03556_ _03402_ _03463_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_17_clk clknet_5_7__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
XFILLER_34_961 VPWR VGND sg13g2_decap_8
X_09342_ VPWR _03494_ _03493_ VGND sg13g2_inv_1
XFILLER_80_588 VPWR VGND sg13g2_decap_8
XFILLER_21_611 VPWR VGND sg13g2_fill_1
XFILLER_33_471 VPWR VGND sg13g2_decap_8
X_09273_ _03427_ _03420_ _03425_ VPWR VGND sg13g2_nand2_1
XFILLER_21_655 VPWR VGND sg13g2_decap_8
XFILLER_32_28 VPWR VGND sg13g2_decap_8
X_08224_ _01371_ _02477_ _02478_ VPWR VGND sg13g2_nand2_1
XFILLER_21_666 VPWR VGND sg13g2_decap_8
XFILLER_119_565 VPWR VGND sg13g2_fill_2
XFILLER_107_705 VPWR VGND sg13g2_decap_4
X_08155_ _02415_ net1659 fp16_sum_pipe.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_20_187 VPWR VGND sg13g2_decap_4
XFILLER_107_738 VPWR VGND sg13g2_decap_8
X_08086_ _02248_ _02351_ _02352_ VPWR VGND sg13g2_nor2_1
XFILLER_115_760 VPWR VGND sg13g2_decap_8
XFILLER_114_270 VPWR VGND sg13g2_decap_8
XFILLER_88_644 VPWR VGND sg13g2_fill_1
XFILLER_0_526 VPWR VGND sg13g2_decap_8
XFILLER_103_988 VPWR VGND sg13g2_decap_8
XFILLER_102_454 VPWR VGND sg13g2_fill_2
XFILLER_87_132 VPWR VGND sg13g2_decap_8
XFILLER_56_530 VPWR VGND sg13g2_decap_8
X_07939_ fp16_sum_pipe.exp_mant_logic0.b\[8\] fp16_sum_pipe.exp_mant_logic0.a\[8\]
+ _02214_ VPWR VGND sg13g2_xor2_1
XFILLER_28_221 VPWR VGND sg13g2_fill_1
XFILLER_28_232 VPWR VGND sg13g2_decap_8
XFILLER_113_42 VPWR VGND sg13g2_decap_8
XFILLER_56_574 VPWR VGND sg13g2_decap_8
XFILLER_16_405 VPWR VGND sg13g2_decap_4
X_10950_ VGND VPWR _04955_ _04864_ _04956_ _04863_ sg13g2_a21oi_1
X_09609_ VPWR _03726_ _03725_ VGND sg13g2_inv_1
XFILLER_44_758 VPWR VGND sg13g2_decap_8
XFILLER_28_287 VPWR VGND sg13g2_fill_2
X_10881_ net1772 _04886_ _04891_ _04892_ VPWR VGND sg13g2_nor3_1
X_12620_ _06436_ _06421_ _05342_ VPWR VGND sg13g2_nand2_1
XFILLER_73_68 VPWR VGND sg13g2_decap_8
XFILLER_71_566 VPWR VGND sg13g2_decap_8
XFILLER_71_544 VPWR VGND sg13g2_decap_8
XFILLER_43_268 VPWR VGND sg13g2_decap_8
XFILLER_43_235 VPWR VGND sg13g2_fill_1
XFILLER_71_599 VPWR VGND sg13g2_decap_4
XFILLER_40_931 VPWR VGND sg13g2_decap_8
XFILLER_25_994 VPWR VGND sg13g2_decap_8
X_12551_ fpdiv.reg_b_out\[15\] fpdiv.reg_a_out\[15\] _06368_ VPWR VGND sg13g2_xor2_1
X_12482_ VGND VPWR _06319_ net1872 _00962_ _06320_ sg13g2_a21oi_1
X_11502_ VPWR _05407_ _05406_ VGND sg13g2_inv_1
XFILLER_125_0 VPWR VGND sg13g2_decap_8
X_11433_ VPWR _05365_ fpdiv.reg_a_out\[10\] VGND sg13g2_inv_1
X_14221_ _00022_ VGND VPWR _00772_ sipo.shift_reg\[2\] clknet_leaf_21_clk sg13g2_dfrbpq_1
XFILLER_8_648 VPWR VGND sg13g2_fill_2
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_11_198 VPWR VGND sg13g2_decap_8
X_14152_ VPWR _00703_ net131 VGND sg13g2_inv_1
XFILLER_125_524 VPWR VGND sg13g2_fill_1
X_11364_ _05314_ _05315_ _05313_ _05316_ VPWR VGND sg13g2_nand3_1
XFILLER_4_832 VPWR VGND sg13g2_decap_8
XFILLER_125_579 VPWR VGND sg13g2_fill_2
X_14083_ VPWR _00634_ net138 VGND sg13g2_inv_1
XFILLER_98_419 VPWR VGND sg13g2_decap_8
X_11295_ _05254_ VPWR _01083_ VGND net1813 _02797_ sg13g2_o21ai_1
X_13103_ _06861_ VPWR _06862_ VGND _06771_ _06801_ sg13g2_o21ai_1
X_10315_ _04375_ net1912 fp16_res_pipe.x2\[8\] VPWR VGND sg13g2_nand2_1
X_13034_ _06802_ _06792_ _06801_ VPWR VGND sg13g2_nand2_2
X_10246_ _04318_ _04317_ net1636 VPWR VGND sg13g2_nand2_1
XFILLER_121_763 VPWR VGND sg13g2_decap_8
XFILLER_120_273 VPWR VGND sg13g2_decap_8
XFILLER_94_614 VPWR VGND sg13g2_decap_8
XFILLER_78_154 VPWR VGND sg13g2_decap_8
X_10177_ VGND VPWR fp16_res_pipe.exp_mant_logic0.a\[2\] net1642 _04256_ _04255_ sg13g2_a21oi_1
XFILLER_94_658 VPWR VGND sg13g2_decap_8
XFILLER_93_124 VPWR VGND sg13g2_fill_2
XFILLER_66_349 VPWR VGND sg13g2_decap_8
XFILLER_14_7 VPWR VGND sg13g2_decap_8
XFILLER_93_168 VPWR VGND sg13g2_decap_4
XFILLER_75_883 VPWR VGND sg13g2_fill_1
XFILLER_62_500 VPWR VGND sg13g2_decap_8
XFILLER_47_552 VPWR VGND sg13g2_decap_8
XFILLER_35_714 VPWR VGND sg13g2_decap_8
XFILLER_35_703 VPWR VGND sg13g2_fill_1
X_13936_ VPWR _00487_ net12 VGND sg13g2_inv_1
XFILLER_62_511 VPWR VGND sg13g2_fill_1
XFILLER_47_596 VPWR VGND sg13g2_fill_2
XFILLER_62_566 VPWR VGND sg13g2_fill_1
X_13867_ VPWR _00418_ net51 VGND sg13g2_inv_1
X_13798_ VPWR _00349_ net73 VGND sg13g2_inv_1
X_12818_ _06600_ VPWR _06601_ VGND net1960 _06598_ sg13g2_o21ai_1
XFILLER_34_279 VPWR VGND sg13g2_decap_8
XFILLER_16_994 VPWR VGND sg13g2_decap_8
X_12749_ fpmul.reg_b_out\[8\] fp16_res_pipe.x2\[8\] net1955 _00918_ VPWR VGND sg13g2_mux2_1
XFILLER_31_942 VPWR VGND sg13g2_decap_8
X_14419_ _00220_ VGND VPWR _00958_ fpmul.seg_reg0.q\[4\] clknet_leaf_78_clk sg13g2_dfrbpq_1
XFILLER_8_63 VPWR VGND sg13g2_decap_8
XFILLER_116_535 VPWR VGND sg13g2_decap_8
XFILLER_7_692 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_6_clk clknet_5_5__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_6_191 VPWR VGND sg13g2_fill_1
X_08911_ _03013_ _02973_ _02998_ _03098_ VPWR VGND sg13g2_nor3_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_98_953 VPWR VGND sg13g2_decap_8
XFILLER_97_441 VPWR VGND sg13g2_decap_8
XFILLER_69_143 VPWR VGND sg13g2_decap_4
X_09891_ fp16_res_pipe.reg1en.q\[0\] _03988_ VPWR VGND sg13g2_inv_4
X_08842_ acc_sub.add_renorm0.mantisa\[11\] acc_sub.add_renorm0.mantisa\[2\] _03029_
+ VPWR VGND sg13g2_nor2_1
XFILLER_112_796 VPWR VGND sg13g2_decap_8
XFILLER_111_273 VPWR VGND sg13g2_decap_4
XFILLER_111_240 VPWR VGND sg13g2_decap_8
XFILLER_97_463 VPWR VGND sg13g2_fill_1
XFILLER_69_165 VPWR VGND sg13g2_decap_8
XFILLER_57_327 VPWR VGND sg13g2_decap_8
XFILLER_111_295 VPWR VGND sg13g2_decap_8
XFILLER_111_284 VPWR VGND sg13g2_fill_1
XFILLER_100_958 VPWR VGND sg13g2_decap_8
X_08773_ _02962_ acc\[1\] net1896 VPWR VGND sg13g2_nand2_1
X_07724_ _01423_ _02029_ _02030_ VPWR VGND sg13g2_nand2_1
XFILLER_84_157 VPWR VGND sg13g2_fill_1
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_65_360 VPWR VGND sg13g2_fill_2
XFILLER_53_533 VPWR VGND sg13g2_decap_8
XFILLER_14_909 VPWR VGND sg13g2_decap_8
XFILLER_26_758 VPWR VGND sg13g2_fill_1
X_07586_ _01900_ _01797_ _01899_ VPWR VGND sg13g2_xnor2_1
XFILLER_43_49 VPWR VGND sg13g2_decap_8
X_09325_ _03478_ fp16_res_pipe.op_sign_logic0.mantisa_a\[9\] fp16_res_pipe.op_sign_logic0.mantisa_b\[9\]
+ VPWR VGND sg13g2_nand2_1
X_09256_ fp16_res_pipe.op_sign_logic0.mantisa_a\[0\] _03409_ _03410_ VPWR VGND sg13g2_nor2_1
XFILLER_22_975 VPWR VGND sg13g2_decap_8
X_08207_ VPWR _02463_ fp16_sum_pipe.exp_mant_logic0.b\[14\] VGND sg13g2_inv_1
X_09187_ _03348_ acc_sub.x2\[5\] net1905 VPWR VGND sg13g2_nand2_1
XFILLER_5_607 VPWR VGND sg13g2_decap_8
XFILLER_119_384 VPWR VGND sg13g2_decap_8
X_08138_ _02399_ net1691 fp16_sum_pipe.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_122_505 VPWR VGND sg13g2_decap_4
X_08069_ _02335_ _02334_ net1652 VPWR VGND sg13g2_nand2_1
Xplace1870 fpmul.reg1en.q\[0\] net1870 VPWR VGND sg13g2_buf_2
Xplace1881 net1880 net1881 VPWR VGND sg13g2_buf_1
X_10100_ _03605_ _04175_ _04184_ VPWR VGND sg13g2_nor2_1
Xplace1892 net1891 net1892 VPWR VGND sg13g2_buf_2
XFILLER_88_441 VPWR VGND sg13g2_decap_4
XFILLER_0_323 VPWR VGND sg13g2_decap_8
XFILLER_1_857 VPWR VGND sg13g2_decap_8
X_10031_ _04118_ _04021_ _04119_ VPWR VGND sg13g2_xor2_1
XFILLER_103_796 VPWR VGND sg13g2_decap_4
XFILLER_103_785 VPWR VGND sg13g2_fill_1
XFILLER_102_262 VPWR VGND sg13g2_decap_4
XFILLER_102_240 VPWR VGND sg13g2_decap_8
XFILLER_89_986 VPWR VGND sg13g2_decap_8
XFILLER_88_463 VPWR VGND sg13g2_decap_8
XFILLER_76_625 VPWR VGND sg13g2_decap_8
XFILLER_48_316 VPWR VGND sg13g2_fill_2
XFILLER_124_63 VPWR VGND sg13g2_decap_8
Xclkbuf_5_26__f_clk clknet_4_13_0_clk clknet_5_26__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_76_669 VPWR VGND sg13g2_decap_4
XFILLER_64_809 VPWR VGND sg13g2_fill_1
XFILLER_84_56 VPWR VGND sg13g2_fill_1
X_14770_ _00571_ VGND VPWR _01294_ acc_sum.exp_mant_logic0.b\[15\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_13721_ VPWR _00272_ net139 VGND sg13g2_inv_1
XFILLER_95_1013 VPWR VGND sg13g2_fill_1
XFILLER_95_1002 VPWR VGND sg13g2_decap_8
XFILLER_72_820 VPWR VGND sg13g2_decap_8
X_11982_ VPWR _05836_ _05835_ VGND sg13g2_inv_1
XFILLER_44_522 VPWR VGND sg13g2_fill_2
X_10933_ VPWR _04940_ fp16_res_pipe.y\[9\] VGND sg13g2_inv_1
XFILLER_32_706 VPWR VGND sg13g2_fill_2
XFILLER_71_374 VPWR VGND sg13g2_fill_1
XFILLER_71_363 VPWR VGND sg13g2_decap_8
X_13652_ VPWR _00203_ net108 VGND sg13g2_inv_1
X_10864_ net1825 fp16_res_pipe.add_renorm0.exp\[5\] _04876_ VPWR VGND sg13g2_nor2_1
X_13583_ VPWR _00134_ net118 VGND sg13g2_inv_1
X_12603_ _06402_ _06397_ _06419_ VPWR VGND sg13g2_xor2_1
X_10795_ fp16_res_pipe.add_renorm0.exp\[2\] _04775_ _04807_ VPWR VGND sg13g2_nor2_1
X_12534_ _06353_ acc_sub.x2\[0\] net1957 VPWR VGND sg13g2_nand2_1
XFILLER_9_913 VPWR VGND sg13g2_decap_8
XFILLER_13_975 VPWR VGND sg13g2_decap_8
XFILLER_40_794 VPWR VGND sg13g2_fill_1
X_12465_ _06307_ _06306_ _06146_ VPWR VGND sg13g2_nand2_1
XFILLER_126_855 VPWR VGND sg13g2_decap_8
X_14204_ VPWR _00755_ net103 VGND sg13g2_inv_1
X_11416_ _05354_ VPWR _01062_ VGND _05353_ net1706 sg13g2_o21ai_1
X_12396_ VGND VPWR _06224_ _06240_ _06242_ _06241_ sg13g2_a21oi_1
X_14135_ VPWR _00686_ net114 VGND sg13g2_inv_1
X_11347_ _05300_ _05297_ _05298_ _05299_ VPWR VGND sg13g2_and3_1
XFILLER_113_538 VPWR VGND sg13g2_decap_8
XFILLER_3_161 VPWR VGND sg13g2_decap_8
X_14066_ VPWR _00617_ net94 VGND sg13g2_inv_1
X_11278_ net1635 VPWR _05240_ VGND _05236_ _05239_ sg13g2_o21ai_1
XFILLER_79_474 VPWR VGND sg13g2_decap_8
X_13017_ _06785_ _06304_ net1853 VPWR VGND sg13g2_nand2_1
X_10229_ _04302_ net1829 VPWR VGND sg13g2_inv_2
XFILLER_95_967 VPWR VGND sg13g2_decap_8
XFILLER_67_658 VPWR VGND sg13g2_decap_4
XFILLER_66_124 VPWR VGND sg13g2_decap_8
XFILLER_39_327 VPWR VGND sg13g2_decap_8
XFILLER_67_669 VPWR VGND sg13g2_decap_8
X_14968_ _00769_ VGND VPWR _01488_ acc_sub.seg_reg1.q\[20\] clknet_leaf_43_clk sg13g2_dfrbpq_1
XFILLER_35_511 VPWR VGND sg13g2_decap_8
X_14899_ _00700_ VGND VPWR _01419_ acc_sub.op_sign_logic0.mantisa_b\[9\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_2
XFILLER_63_875 VPWR VGND sg13g2_decap_8
X_13919_ VPWR _00470_ net5 VGND sg13g2_inv_1
X_07440_ VPWR _01770_ fpdiv.divider0.divisor_reg\[6\] VGND sg13g2_inv_1
XFILLER_90_661 VPWR VGND sg13g2_decap_4
X_07371_ acc_sub.add_renorm0.exp\[0\] acc_sub.seg_reg0.q\[22\] net1797 _01468_ VPWR
+ VGND sg13g2_mux2_1
X_09110_ net1786 VPWR _03292_ VGND _03291_ _03231_ sg13g2_o21ai_1
XFILLER_88_0 VPWR VGND sg13g2_decap_8
XFILLER_50_569 VPWR VGND sg13g2_decap_4
XFILLER_31_750 VPWR VGND sg13g2_fill_2
X_09041_ _03080_ _03226_ _03227_ VPWR VGND sg13g2_nor2b_1
XFILLER_117_844 VPWR VGND sg13g2_decap_8
XFILLER_104_527 VPWR VGND sg13g2_fill_2
XFILLER_104_549 VPWR VGND sg13g2_decap_8
X_09943_ _04019_ VPWR _04039_ VGND _04033_ _04038_ sg13g2_o21ai_1
XFILLER_112_560 VPWR VGND sg13g2_fill_1
X_09874_ net1820 acc_sum.y\[4\] _03980_ VPWR VGND sg13g2_nor2_1
XFILLER_100_700 VPWR VGND sg13g2_fill_1
X_08825_ VGND VPWR _03010_ _02996_ _03012_ _03011_ sg13g2_a21oi_1
XFILLER_100_744 VPWR VGND sg13g2_fill_2
XFILLER_86_945 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_decap_8
XFILLER_79_1008 VPWR VGND sg13g2_decap_4
XFILLER_73_617 VPWR VGND sg13g2_decap_8
XFILLER_45_308 VPWR VGND sg13g2_decap_8
XFILLER_39_861 VPWR VGND sg13g2_decap_8
X_08756_ _02950_ VPWR _01318_ VGND net1898 _02949_ sg13g2_o21ai_1
XFILLER_45_319 VPWR VGND sg13g2_fill_1
X_07707_ _01745_ _01977_ _02014_ VPWR VGND sg13g2_nor2_1
X_08687_ net1668 VPWR _02902_ VGND _02748_ _02901_ sg13g2_o21ai_1
XFILLER_72_138 VPWR VGND sg13g2_decap_8
XFILLER_26_533 VPWR VGND sg13g2_fill_1
XFILLER_26_566 VPWR VGND sg13g2_fill_2
XFILLER_26_588 VPWR VGND sg13g2_decap_4
XFILLER_110_21 VPWR VGND sg13g2_decap_8
X_07569_ _01882_ VPWR _01883_ VGND acc_sub.exp_mant_logic0.a\[8\] _01825_ sg13g2_o21ai_1
XFILLER_41_547 VPWR VGND sg13g2_decap_4
X_09308_ _03460_ VPWR _03461_ VGND _03412_ _03414_ sg13g2_o21ai_1
XFILLER_10_912 VPWR VGND sg13g2_decap_8
X_10580_ _04603_ acc_sub.x2\[9\] net1925 VPWR VGND sg13g2_nand2_1
XFILLER_6_927 VPWR VGND sg13g2_decap_8
X_09239_ fp16_res_pipe.op_sign_logic0.mantisa_a\[5\] _03392_ _03393_ VPWR VGND sg13g2_nor2_1
XFILLER_119_63 VPWR VGND sg13g2_decap_8
X_12250_ _06096_ _06095_ _05961_ VPWR VGND sg13g2_nand2b_1
XFILLER_5_415 VPWR VGND sg13g2_fill_2
XFILLER_10_989 VPWR VGND sg13g2_decap_8
XFILLER_79_23 VPWR VGND sg13g2_decap_8
X_11201_ _05168_ net1809 net1655 net1810 _05124_ VPWR VGND sg13g2_a22oi_1
X_12181_ _05998_ _05993_ _06027_ VPWR VGND sg13g2_and2_1
XFILLER_122_324 VPWR VGND sg13g2_fill_2
X_11132_ _05086_ _05048_ _05102_ VPWR VGND sg13g2_nor2_1
XFILLER_123_869 VPWR VGND sg13g2_decap_8
XFILLER_96_709 VPWR VGND sg13g2_decap_8
XFILLER_95_219 VPWR VGND sg13g2_fill_2
X_11063_ VPWR VGND _05039_ _05040_ _05036_ acc_sum.exp_mant_logic0.a\[14\] _05041_
+ _03329_ sg13g2_a221oi_1
XFILLER_62_1012 VPWR VGND sg13g2_fill_2
XFILLER_49_614 VPWR VGND sg13g2_decap_4
XFILLER_103_582 VPWR VGND sg13g2_decap_8
XFILLER_89_794 VPWR VGND sg13g2_decap_8
XFILLER_88_293 VPWR VGND sg13g2_decap_4
XFILLER_49_658 VPWR VGND sg13g2_fill_1
X_10014_ _04102_ _04008_ _04101_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_175 VPWR VGND sg13g2_decap_8
X_14822_ _00623_ VGND VPWR _01346_ acc_sum.add_renorm0.mantisa\[11\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_2
XFILLER_95_99 VPWR VGND sg13g2_fill_1
XFILLER_95_77 VPWR VGND sg13g2_decap_8
XFILLER_91_414 VPWR VGND sg13g2_fill_1
XFILLER_57_691 VPWR VGND sg13g2_fill_2
X_14753_ _00554_ VGND VPWR net1813 acc_sum.reg2en.q\[0\] clknet_leaf_32_clk sg13g2_dfrbpq_2
X_11965_ _05820_ VPWR _00979_ VGND net1883 _05819_ sg13g2_o21ai_1
XFILLER_72_661 VPWR VGND sg13g2_fill_2
X_13704_ VPWR _00255_ net65 VGND sg13g2_inv_1
X_14684_ _00485_ VGND VPWR _01212_ fp16_res_pipe.op_sign_logic0.mantisa_a\[10\] clknet_leaf_139_clk
+ sg13g2_dfrbpq_1
X_10916_ _04924_ _04862_ _04925_ VPWR VGND sg13g2_nor2b_1
XFILLER_71_171 VPWR VGND sg13g2_fill_2
X_13635_ VPWR _00186_ net61 VGND sg13g2_inv_1
X_11896_ fpmul.seg_reg0.q\[52\] fpmul.reg_a_out\[13\] net1878 _01006_ VPWR VGND sg13g2_mux2_1
XFILLER_44_70 VPWR VGND sg13g2_decap_8
XFILLER_60_878 VPWR VGND sg13g2_fill_2
X_10847_ net1825 _03576_ _04859_ VPWR VGND sg13g2_nor2_1
X_13566_ VPWR _00117_ net33 VGND sg13g2_inv_1
XFILLER_9_732 VPWR VGND sg13g2_decap_4
XFILLER_13_772 VPWR VGND sg13g2_decap_8
X_10778_ _04790_ _04786_ fp16_res_pipe.add_renorm0.exp\[5\] VPWR VGND sg13g2_nand2_1
X_13497_ VPWR _00048_ net33 VGND sg13g2_inv_1
X_12517_ fpmul.reg_a_out\[8\] net1955 _06344_ VPWR VGND sg13g2_nor2_1
XFILLER_40_591 VPWR VGND sg13g2_decap_8
X_12448_ _00969_ _06292_ _06293_ VPWR VGND sg13g2_nand2_1
XFILLER_126_663 VPWR VGND sg13g2_fill_1
XFILLER_125_140 VPWR VGND sg13g2_decap_8
XFILLER_99_503 VPWR VGND sg13g2_decap_8
XFILLER_114_825 VPWR VGND sg13g2_decap_8
XFILLER_113_302 VPWR VGND sg13g2_fill_2
XFILLER_99_536 VPWR VGND sg13g2_decap_4
X_12379_ _06225_ net1858 fpmul.reg_b_out\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_5_42 VPWR VGND sg13g2_decap_8
XFILLER_99_547 VPWR VGND sg13g2_fill_2
X_14118_ VPWR _00669_ net46 VGND sg13g2_inv_1
XFILLER_86_219 VPWR VGND sg13g2_decap_4
XFILLER_67_400 VPWR VGND sg13g2_decap_4
X_14049_ VPWR _00600_ net23 VGND sg13g2_inv_1
XFILLER_68_945 VPWR VGND sg13g2_fill_1
X_08610_ acc_sum.op_sign_logic0.mantisa_a\[7\] acc_sum.op_sign_logic0.mantisa_b\[7\]
+ net1740 _02833_ VPWR VGND sg13g2_nand3_1
XFILLER_83_904 VPWR VGND sg13g2_decap_8
XFILLER_28_809 VPWR VGND sg13g2_decap_8
X_09590_ _03704_ _03706_ _03701_ _03707_ VPWR VGND sg13g2_nand3_1
XFILLER_94_263 VPWR VGND sg13g2_fill_1
X_08541_ VPWR _02765_ _02764_ VGND sg13g2_inv_1
XFILLER_70_609 VPWR VGND sg13g2_decap_4
XFILLER_47_190 VPWR VGND sg13g2_decap_8
XFILLER_36_842 VPWR VGND sg13g2_fill_2
X_08472_ _02703_ net1647 _02702_ VPWR VGND sg13g2_nand2_1
XFILLER_51_812 VPWR VGND sg13g2_decap_8
XFILLER_50_300 VPWR VGND sg13g2_fill_1
XFILLER_36_875 VPWR VGND sg13g2_decap_4
X_07423_ VPWR _01758_ _01756_ VGND sg13g2_inv_1
XFILLER_63_694 VPWR VGND sg13g2_fill_1
XFILLER_62_171 VPWR VGND sg13g2_fill_2
X_07354_ _01712_ net1797 acc_sub.seg_reg0.q\[28\] VPWR VGND sg13g2_nand2_1
XFILLER_10_208 VPWR VGND sg13g2_decap_8
X_07285_ VGND VPWR _01652_ _01507_ _01653_ _01635_ sg13g2_a21oi_1
X_09024_ _03183_ _03209_ _03210_ VPWR VGND sg13g2_nor2_1
XFILLER_117_630 VPWR VGND sg13g2_fill_2
XFILLER_40_28 VPWR VGND sg13g2_decap_8
XFILLER_116_173 VPWR VGND sg13g2_decap_8
XFILLER_120_806 VPWR VGND sg13g2_decap_8
X_09926_ _04023_ _04022_ fp16_res_pipe.exp_mant_logic0.a\[9\] VPWR VGND sg13g2_nand2_1
X_09857_ VPWR _03966_ acc_sum.y\[7\] VGND sg13g2_inv_1
X_08808_ _02995_ _02994_ VPWR VGND sg13g2_inv_2
X_09788_ VPWR _03902_ _03819_ VGND sg13g2_inv_1
XFILLER_86_786 VPWR VGND sg13g2_decap_8
XFILLER_73_403 VPWR VGND sg13g2_decap_4
XFILLER_46_628 VPWR VGND sg13g2_decap_4
XFILLER_45_105 VPWR VGND sg13g2_decap_8
X_08739_ VPWR _02939_ acc_sum.exp_mant_logic0.a\[12\] VGND sg13g2_inv_1
XFILLER_27_853 VPWR VGND sg13g2_decap_8
XFILLER_121_42 VPWR VGND sg13g2_decap_8
X_11750_ _05653_ VPWR _05654_ VGND net1839 fp16_sum_pipe.add_renorm0.exp\[6\] sg13g2_o21ai_1
XFILLER_26_374 VPWR VGND sg13g2_decap_8
XFILLER_27_897 VPWR VGND sg13g2_decap_8
X_10701_ _04713_ VPWR _04714_ VGND net1826 _04656_ sg13g2_o21ai_1
XFILLER_14_536 VPWR VGND sg13g2_decap_4
XFILLER_26_385 VPWR VGND sg13g2_fill_2
XFILLER_14_569 VPWR VGND sg13g2_fill_2
X_13420_ _07089_ net1720 instr\[7\] VPWR VGND sg13g2_nand2_1
X_10632_ fp16_res_pipe.add_renorm0.mantisa\[4\] fp16_res_pipe.add_renorm0.mantisa\[3\]
+ fp16_res_pipe.add_renorm0.mantisa\[5\] _04645_ VPWR VGND fp16_res_pipe.add_renorm0.mantisa\[2\]
+ sg13g2_nand4_1
XFILLER_22_580 VPWR VGND sg13g2_fill_2
X_13351_ _07049_ VPWR _00823_ VGND _07003_ net1724 sg13g2_o21ai_1
XFILLER_10_753 VPWR VGND sg13g2_fill_1
XFILLER_14_84 VPWR VGND sg13g2_fill_1
X_10563_ _04594_ fp16_sum_pipe.seg_reg0.q\[23\] net1845 VPWR VGND sg13g2_nand2_1
X_12302_ _06059_ _06147_ _06148_ VPWR VGND sg13g2_nor2_1
XFILLER_6_735 VPWR VGND sg13g2_fill_1
XFILLER_5_201 VPWR VGND sg13g2_fill_1
X_13282_ VGND VPWR net1676 _06997_ _00841_ _06998_ sg13g2_a21oi_1
XFILLER_5_223 VPWR VGND sg13g2_fill_2
X_10494_ VGND VPWR _04538_ _04408_ _04539_ _04405_ sg13g2_a21oi_1
XFILLER_108_696 VPWR VGND sg13g2_decap_8
XFILLER_107_140 VPWR VGND sg13g2_decap_8
X_12233_ _06079_ net1856 net1867 VPWR VGND sg13g2_nand2_1
XFILLER_5_256 VPWR VGND sg13g2_fill_1
X_12164_ _06007_ _05983_ _06005_ _06010_ VPWR VGND sg13g2_nand3_1
XFILLER_122_154 VPWR VGND sg13g2_decap_8
XFILLER_111_817 VPWR VGND sg13g2_decap_8
XFILLER_96_506 VPWR VGND sg13g2_decap_4
X_11115_ VPWR _05085_ _05084_ VGND sg13g2_inv_1
X_12095_ VPWR _05941_ _05897_ VGND sg13g2_inv_1
XFILLER_110_316 VPWR VGND sg13g2_decap_8
X_11046_ _05018_ _05024_ _05025_ VPWR VGND sg13g2_nor2_1
XFILLER_2_996 VPWR VGND sg13g2_decap_8
XFILLER_77_775 VPWR VGND sg13g2_fill_1
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_91_200 VPWR VGND sg13g2_decap_8
XFILLER_65_959 VPWR VGND sg13g2_decap_8
XFILLER_49_477 VPWR VGND sg13g2_fill_1
XFILLER_36_105 VPWR VGND sg13g2_decap_8
XFILLER_92_767 VPWR VGND sg13g2_decap_8
X_14805_ _00606_ VGND VPWR _01329_ acc_sum.add_renorm0.exp\[2\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_18_842 VPWR VGND sg13g2_fill_2
X_12997_ VPWR _06765_ _06764_ VGND sg13g2_inv_1
XFILLER_55_80 VPWR VGND sg13g2_decap_8
X_14736_ _00537_ VGND VPWR _01264_ fp16_res_pipe.add_renorm0.exp\[7\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_1
XFILLER_18_864 VPWR VGND sg13g2_fill_1
XFILLER_91_299 VPWR VGND sg13g2_decap_4
XFILLER_73_992 VPWR VGND sg13g2_fill_1
X_11948_ VPWR _05809_ fpmul.seg_reg0.q\[30\] VGND sg13g2_inv_1
X_11879_ _05768_ fpdiv.divider0.counter\[1\] fpdiv.divider0.counter\[0\] VPWR VGND
+ sg13g2_nand2_1
XFILLER_60_664 VPWR VGND sg13g2_decap_8
XFILLER_60_653 VPWR VGND sg13g2_fill_1
X_14667_ _00468_ VGND VPWR _01195_ fp16_res_pipe.op_sign_logic0.mantisa_b\[4\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_2
X_13618_ VPWR _00169_ net61 VGND sg13g2_inv_1
X_14598_ _00399_ VGND VPWR _01130_ fp16_res_pipe.y\[9\] clknet_leaf_129_clk sg13g2_dfrbpq_1
XFILLER_32_388 VPWR VGND sg13g2_decap_8
XFILLER_32_399 VPWR VGND sg13g2_fill_2
X_13549_ VPWR _00100_ net88 VGND sg13g2_inv_1
XFILLER_9_562 VPWR VGND sg13g2_decap_8
XFILLER_118_438 VPWR VGND sg13g2_decap_4
XFILLER_114_622 VPWR VGND sg13g2_fill_1
XFILLER_114_600 VPWR VGND sg13g2_decap_8
XFILLER_114_688 VPWR VGND sg13g2_decap_8
XFILLER_102_817 VPWR VGND sg13g2_fill_1
XFILLER_101_305 VPWR VGND sg13g2_fill_2
XFILLER_87_506 VPWR VGND sg13g2_decap_8
XFILLER_101_338 VPWR VGND sg13g2_decap_8
X_09711_ _03826_ _03785_ _03827_ VPWR VGND sg13g2_nor2_1
X_07972_ _02244_ _02245_ VPWR VGND sg13g2_inv_4
XFILLER_110_850 VPWR VGND sg13g2_decap_8
XFILLER_28_606 VPWR VGND sg13g2_decap_8
X_09642_ _03759_ _03717_ _03758_ VPWR VGND sg13g2_nand2b_1
XFILLER_55_425 VPWR VGND sg13g2_decap_4
XFILLER_27_105 VPWR VGND sg13g2_decap_8
X_09573_ _03690_ net1806 acc_sum.add_renorm0.mantisa\[7\] VPWR VGND sg13g2_nand2_1
X_08524_ acc_sum.op_sign_logic0.mantisa_a\[2\] _02747_ _02748_ VPWR VGND sg13g2_nor2_2
XFILLER_35_28 VPWR VGND sg13g2_decap_8
XFILLER_70_428 VPWR VGND sg13g2_decap_8
XFILLER_42_119 VPWR VGND sg13g2_decap_8
XFILLER_36_683 VPWR VGND sg13g2_decap_8
XFILLER_35_182 VPWR VGND sg13g2_fill_1
XFILLER_24_845 VPWR VGND sg13g2_decap_4
X_08455_ _02688_ VPWR _01357_ VGND net1705 _02686_ sg13g2_o21ai_1
XFILLER_51_664 VPWR VGND sg13g2_fill_1
XFILLER_51_642 VPWR VGND sg13g2_fill_2
XFILLER_23_344 VPWR VGND sg13g2_fill_2
X_07406_ _01746_ net1894 acc\[4\] VPWR VGND sg13g2_nand2_1
X_08386_ _02624_ _07113_ _02623_ VPWR VGND sg13g2_nand2_1
XFILLER_50_185 VPWR VGND sg13g2_fill_2
XFILLER_23_377 VPWR VGND sg13g2_decap_8
X_07337_ _01699_ _01697_ _01698_ acc_sub.add_renorm0.mantisa\[2\] net1784 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_51_49 VPWR VGND sg13g2_decap_8
XFILLER_109_416 VPWR VGND sg13g2_decap_4
XFILLER_118_950 VPWR VGND sg13g2_decap_8
X_07268_ _01622_ _01637_ _01621_ _01486_ VPWR VGND sg13g2_nand3_1
XFILLER_124_408 VPWR VGND sg13g2_fill_2
X_07199_ VPWR _01571_ _01570_ VGND sg13g2_inv_1
XFILLER_117_460 VPWR VGND sg13g2_decap_8
X_09007_ VPWR _03193_ _03149_ VGND sg13g2_inv_1
XFILLER_105_611 VPWR VGND sg13g2_decap_8
XFILLER_105_644 VPWR VGND sg13g2_fill_1
XFILLER_3_749 VPWR VGND sg13g2_decap_8
XFILLER_120_614 VPWR VGND sg13g2_decap_4
XFILLER_78_528 VPWR VGND sg13g2_decap_4
XFILLER_116_75 VPWR VGND sg13g2_decap_8
XFILLER_105_699 VPWR VGND sg13g2_fill_1
XFILLER_120_658 VPWR VGND sg13g2_decap_8
XFILLER_58_230 VPWR VGND sg13g2_decap_8
X_09909_ fp16_res_pipe.exp_mant_logic0.a\[11\] _04005_ _04006_ VPWR VGND sg13g2_nor2_1
X_12920_ VGND VPWR net1936 add_result\[4\] _06694_ net1950 sg13g2_a21oi_1
XFILLER_46_425 VPWR VGND sg13g2_fill_1
XFILLER_46_414 VPWR VGND sg13g2_decap_8
XFILLER_73_244 VPWR VGND sg13g2_decap_4
X_12851_ _06631_ _06630_ _06629_ VPWR VGND sg13g2_nand2b_1
XFILLER_18_149 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
X_11802_ _01025_ _05702_ _05703_ VPWR VGND sg13g2_nand2_1
XFILLER_109_1012 VPWR VGND sg13g2_fill_2
XFILLER_92_67 VPWR VGND sg13g2_fill_2
X_12782_ VPWR _06567_ _06566_ VGND sg13g2_inv_1
XFILLER_55_992 VPWR VGND sg13g2_fill_1
XFILLER_54_491 VPWR VGND sg13g2_fill_2
XFILLER_42_620 VPWR VGND sg13g2_decap_8
XFILLER_70_951 VPWR VGND sg13g2_decap_8
X_14521_ _00322_ VGND VPWR _01057_ fpdiv.reg_a_out\[12\] clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_42_653 VPWR VGND sg13g2_decap_8
XFILLER_14_333 VPWR VGND sg13g2_fill_1
XFILLER_15_889 VPWR VGND sg13g2_decap_8
X_11733_ _05617_ _05488_ _05637_ VPWR VGND sg13g2_nor2_1
X_14452_ _00253_ VGND VPWR _00991_ fpmul.seg_reg0.q\[37\] clknet_leaf_122_clk sg13g2_dfrbpq_1
X_11664_ _05555_ _05563_ _05568_ _05569_ VPWR VGND sg13g2_nor3_1
XFILLER_30_848 VPWR VGND sg13g2_decap_8
X_13403_ _07080_ net1721 instr\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_41_185 VPWR VGND sg13g2_fill_2
X_10615_ VPWR _04628_ fp16_res_pipe.add_renorm0.mantisa\[3\] VGND sg13g2_inv_1
XFILLER_127_224 VPWR VGND sg13g2_decap_8
X_14383_ _00184_ VGND VPWR _00924_ fpmul.reg_b_out\[14\] clknet_leaf_124_clk sg13g2_dfrbpq_1
X_11595_ VGND VPWR _05489_ _05497_ _05500_ net1757 sg13g2_a21oi_1
X_13334_ _07039_ net1726 fp16_res_pipe.x2\[11\] VPWR VGND sg13g2_nand2_1
X_10546_ _04582_ VPWR _01160_ VGND net1846 _04581_ sg13g2_o21ai_1
XFILLER_115_408 VPWR VGND sg13g2_decap_4
X_13265_ VGND VPWR net1679 _06984_ _00845_ _06985_ sg13g2_a21oi_1
X_10477_ VGND VPWR _04515_ _04453_ _04524_ _04452_ sg13g2_a21oi_1
XFILLER_124_942 VPWR VGND sg13g2_decap_8
XFILLER_108_482 VPWR VGND sg13g2_fill_1
X_12216_ _06020_ _06061_ _06056_ _06062_ VPWR VGND sg13g2_nand3_1
XFILLER_44_7 VPWR VGND sg13g2_decap_8
XFILLER_29_1013 VPWR VGND sg13g2_fill_1
XFILLER_123_452 VPWR VGND sg13g2_decap_8
X_13196_ _06932_ net1713 sipo.word\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_110_113 VPWR VGND sg13g2_decap_4
XFILLER_110_102 VPWR VGND sg13g2_fill_2
XFILLER_97_859 VPWR VGND sg13g2_decap_8
XFILLER_69_539 VPWR VGND sg13g2_decap_4
X_12147_ fpmul.reg_a_out\[3\] fpmul.reg_b_out\[6\] net1856 _05993_ VPWR VGND sg13g2_nand3_1
XFILLER_2_793 VPWR VGND sg13g2_decap_8
X_12078_ _05924_ _05921_ _05923_ VPWR VGND sg13g2_nand2_1
XFILLER_38_904 VPWR VGND sg13g2_decap_8
XFILLER_1_292 VPWR VGND sg13g2_decap_8
XFILLER_2_21 VPWR VGND sg13g2_decap_8
X_11029_ acc_sum.exp_mant_logic0.b\[13\] _02937_ _05008_ VPWR VGND sg13g2_nor2_1
XFILLER_64_211 VPWR VGND sg13g2_decap_4
XFILLER_38_959 VPWR VGND sg13g2_decap_8
XFILLER_2_98 VPWR VGND sg13g2_decap_8
XFILLER_92_564 VPWR VGND sg13g2_fill_1
XFILLER_65_789 VPWR VGND sg13g2_decap_8
XFILLER_18_672 VPWR VGND sg13g2_decap_8
XFILLER_64_299 VPWR VGND sg13g2_decap_8
XFILLER_21_804 VPWR VGND sg13g2_decap_8
X_14719_ _00520_ VGND VPWR _01247_ fp16_res_pipe.exp_mant_logic0.a\[6\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
XFILLER_33_642 VPWR VGND sg13g2_fill_1
XFILLER_123_1009 VPWR VGND sg13g2_decap_4
XFILLER_60_472 VPWR VGND sg13g2_fill_2
XFILLER_33_675 VPWR VGND sg13g2_decap_8
X_08240_ _02492_ net1658 _02472_ VPWR VGND sg13g2_nand2_1
XFILLER_32_163 VPWR VGND sg13g2_fill_1
XFILLER_20_336 VPWR VGND sg13g2_decap_8
X_08171_ _02428_ _02429_ _02430_ VPWR VGND sg13g2_nor2b_1
X_07122_ _01495_ acc_sub.op_sign_logic0.add_sub _01494_ VPWR VGND sg13g2_xnor2_1
XFILLER_70_0 VPWR VGND sg13g2_decap_8
XFILLER_119_758 VPWR VGND sg13g2_decap_8
XFILLER_118_224 VPWR VGND sg13g2_decap_8
XFILLER_115_942 VPWR VGND sg13g2_decap_8
XFILLER_114_485 VPWR VGND sg13g2_decap_4
XFILLER_102_625 VPWR VGND sg13g2_fill_2
XFILLER_102_614 VPWR VGND sg13g2_decap_8
XFILLER_101_113 VPWR VGND sg13g2_decap_8
XFILLER_87_336 VPWR VGND sg13g2_decap_8
Xclkbuf_5_7__f_clk clknet_4_3_0_clk clknet_5_7__leaf_clk VPWR VGND sg13g2_buf_8
X_07955_ _02228_ VPWR _02229_ VGND _02217_ _02214_ sg13g2_o21ai_1
XFILLER_96_892 VPWR VGND sg13g2_decap_4
XFILLER_29_948 VPWR VGND sg13g2_decap_8
X_09625_ _03742_ _03696_ _03719_ VPWR VGND sg13g2_xnor2_1
X_07886_ _02170_ net1892 acc_sub.x2\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_44_907 VPWR VGND sg13g2_decap_8
XFILLER_56_789 VPWR VGND sg13g2_fill_1
X_09556_ _03673_ acc_sum.add_renorm0.mantisa\[3\] VPWR VGND sg13g2_inv_2
XFILLER_70_214 VPWR VGND sg13g2_fill_1
XFILLER_55_299 VPWR VGND sg13g2_decap_8
XFILLER_36_480 VPWR VGND sg13g2_decap_8
XFILLER_15_119 VPWR VGND sg13g2_fill_2
XFILLER_24_620 VPWR VGND sg13g2_fill_2
XFILLER_102_66 VPWR VGND sg13g2_decap_8
X_08507_ acc_sum.op_sign_logic0.mantisa_b\[9\] acc_sum.op_sign_logic0.mantisa_a\[9\]
+ _02731_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_940 VPWR VGND sg13g2_decap_4
XFILLER_24_664 VPWR VGND sg13g2_decap_8
X_09487_ _03609_ fp16_res_pipe.exp_mant_logic0.a\[4\] VPWR VGND sg13g2_inv_2
X_08438_ _02672_ fpdiv.divider0.divisor_reg\[8\] fpdiv.divider0.remainder_reg\[8\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_62_59 VPWR VGND sg13g2_fill_2
XFILLER_51_483 VPWR VGND sg13g2_decap_8
XFILLER_24_675 VPWR VGND sg13g2_fill_1
XFILLER_12_848 VPWR VGND sg13g2_decap_8
X_08369_ VPWR _02612_ instr\[0\] VGND sg13g2_inv_1
X_11380_ _01074_ _05329_ _05330_ VPWR VGND sg13g2_nand2_1
X_10400_ _04449_ VPWR _04450_ VGND _04411_ _04448_ sg13g2_o21ai_1
XFILLER_20_892 VPWR VGND sg13g2_decap_8
XFILLER_125_739 VPWR VGND sg13g2_decap_8
X_10331_ _04383_ net1921 fp16_res_pipe.x2\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_124_238 VPWR VGND sg13g2_decap_8
X_13050_ _05863_ _06749_ _06754_ _06818_ VPWR VGND sg13g2_nor3_1
XFILLER_3_546 VPWR VGND sg13g2_decap_8
XFILLER_11_63 VPWR VGND sg13g2_decap_8
X_10262_ _04333_ _04325_ _04332_ VPWR VGND sg13g2_nand2_1
XFILLER_127_63 VPWR VGND sg13g2_decap_8
XFILLER_106_964 VPWR VGND sg13g2_decap_8
X_12001_ fpmul.reg_b_out\[13\] fpmul.reg_a_out\[13\] _05855_ VPWR VGND sg13g2_xor2_1
XFILLER_121_945 VPWR VGND sg13g2_decap_8
XFILLER_120_411 VPWR VGND sg13g2_decap_4
X_10193_ _04270_ VPWR _01201_ VGND net1831 _03368_ sg13g2_o21ai_1
XFILLER_78_358 VPWR VGND sg13g2_decap_8
X_13952_ VPWR _00503_ net98 VGND sg13g2_inv_1
XFILLER_94_829 VPWR VGND sg13g2_decap_8
XFILLER_59_572 VPWR VGND sg13g2_decap_8
XFILLER_19_403 VPWR VGND sg13g2_fill_1
X_12903_ _06678_ VPWR _06679_ VGND net1962 _06676_ sg13g2_o21ai_1
XFILLER_46_211 VPWR VGND sg13g2_decap_8
XFILLER_74_553 VPWR VGND sg13g2_decap_8
XFILLER_62_704 VPWR VGND sg13g2_fill_1
XFILLER_35_918 VPWR VGND sg13g2_decap_8
X_13883_ VPWR _00434_ net48 VGND sg13g2_inv_1
X_12834_ _00017_ net1730 net1701 _06615_ VPWR VGND sg13g2_nand3_1
XFILLER_74_586 VPWR VGND sg13g2_fill_2
XFILLER_46_288 VPWR VGND sg13g2_fill_1
XFILLER_15_620 VPWR VGND sg13g2_fill_2
XFILLER_27_480 VPWR VGND sg13g2_decap_8
X_12765_ _06549_ VPWR _06550_ VGND net1923 _06548_ sg13g2_o21ai_1
X_14504_ _00305_ VGND VPWR _01040_ fpdiv.reg_b_out\[11\] clknet_leaf_91_clk sg13g2_dfrbpq_2
X_11716_ VGND VPWR _05493_ _05596_ _05620_ _05619_ sg13g2_a21oi_1
X_12696_ _06435_ _06437_ _06505_ VPWR VGND sg13g2_nor2_1
XFILLER_42_483 VPWR VGND sg13g2_decap_4
X_14435_ _00236_ VGND VPWR _00974_ fpmul.seg_reg0.q\[20\] clknet_leaf_96_clk sg13g2_dfrbpq_1
X_11647_ _05552_ _05434_ _05465_ _05470_ _05442_ VPWR VGND sg13g2_a22oi_1
X_14366_ _00167_ VGND VPWR _00908_ _00019_ clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_10_380 VPWR VGND sg13g2_decap_8
X_11578_ _05428_ _05482_ _05462_ _05483_ VPWR VGND sg13g2_nor3_2
X_13317_ VPWR _07026_ sipo.word\[15\] VGND sg13g2_inv_1
XFILLER_7_874 VPWR VGND sg13g2_decap_8
XFILLER_6_362 VPWR VGND sg13g2_decap_8
X_10529_ _04569_ net1673 _04418_ VPWR VGND sg13g2_nand2b_1
XFILLER_115_238 VPWR VGND sg13g2_decap_8
X_14297_ _00098_ VGND VPWR _00841_ acc\[7\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_112_901 VPWR VGND sg13g2_decap_8
XFILLER_69_303 VPWR VGND sg13g2_decap_8
X_13179_ VPWR _06920_ sipo.shift_reg\[11\] VGND sg13g2_inv_1
XFILLER_112_978 VPWR VGND sg13g2_decap_8
XFILLER_57_509 VPWR VGND sg13g2_decap_8
X_07740_ _02045_ _02043_ _02044_ VPWR VGND sg13g2_nand2_1
XFILLER_93_840 VPWR VGND sg13g2_decap_8
X_07671_ _01973_ _01978_ _01980_ _01981_ VPWR VGND sg13g2_nor3_1
XFILLER_93_884 VPWR VGND sg13g2_decap_8
XFILLER_80_501 VPWR VGND sg13g2_fill_1
XFILLER_53_715 VPWR VGND sg13g2_decap_8
X_09410_ _03555_ _03361_ fp16_res_pipe.add_renorm0.mantisa\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_19_992 VPWR VGND sg13g2_decap_8
XFILLER_25_417 VPWR VGND sg13g2_decap_8
XFILLER_80_545 VPWR VGND sg13g2_fill_1
XFILLER_52_236 VPWR VGND sg13g2_decap_8
XFILLER_40_409 VPWR VGND sg13g2_decap_8
XFILLER_34_940 VPWR VGND sg13g2_decap_8
X_09341_ VGND VPWR _03492_ _03428_ _03493_ _03395_ sg13g2_a21oi_1
XFILLER_60_291 VPWR VGND sg13g2_decap_8
XFILLER_60_280 VPWR VGND sg13g2_decap_8
XFILLER_21_645 VPWR VGND sg13g2_fill_1
XFILLER_119_511 VPWR VGND sg13g2_decap_8
X_08223_ _02478_ fp16_sum_pipe.exp_mant_logic0.b\[6\] _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[9\]
+ net1777 VPWR VGND sg13g2_a22oi_1
XFILLER_119_544 VPWR VGND sg13g2_decap_8
X_08154_ _02267_ _02396_ _02414_ VPWR VGND sg13g2_nor2_1
XFILLER_20_177 VPWR VGND sg13g2_fill_2
XFILLER_119_588 VPWR VGND sg13g2_fill_2
XFILLER_119_577 VPWR VGND sg13g2_decap_8
X_08085_ _02330_ _02335_ _02350_ _02351_ VPWR VGND sg13g2_nor3_1
XFILLER_0_505 VPWR VGND sg13g2_decap_8
XFILLER_103_967 VPWR VGND sg13g2_decap_8
X_08987_ VGND VPWR _03172_ _03173_ _03171_ _03146_ sg13g2_a21oi_2
Xclkbuf_4_5_0_clk clknet_0_clk clknet_4_5_0_clk VPWR VGND sg13g2_buf_8
XFILLER_29_712 VPWR VGND sg13g2_fill_1
XFILLER_113_21 VPWR VGND sg13g2_decap_8
XFILLER_87_188 VPWR VGND sg13g2_fill_2
XFILLER_69_892 VPWR VGND sg13g2_fill_2
XFILLER_28_200 VPWR VGND sg13g2_decap_8
X_07938_ _02213_ _02207_ _02212_ VPWR VGND sg13g2_nand2_1
X_07869_ _02161_ VPWR _01409_ VGND net1885 _01776_ sg13g2_o21ai_1
XFILLER_113_98 VPWR VGND sg13g2_decap_8
X_09608_ _03724_ VPWR _03725_ VGND net1805 _03619_ sg13g2_o21ai_1
XFILLER_84_895 VPWR VGND sg13g2_fill_2
XFILLER_73_36 VPWR VGND sg13g2_decap_8
XFILLER_44_737 VPWR VGND sg13g2_decap_8
XFILLER_43_214 VPWR VGND sg13g2_decap_8
XFILLER_16_417 VPWR VGND sg13g2_decap_8
X_10880_ VGND VPWR _04890_ _04831_ _04891_ _04742_ sg13g2_a21oi_1
XFILLER_52_770 VPWR VGND sg13g2_fill_1
XFILLER_12_601 VPWR VGND sg13g2_decap_8
XFILLER_24_450 VPWR VGND sg13g2_decap_8
XFILLER_25_973 VPWR VGND sg13g2_decap_8
X_12481_ net1872 fpmul.seg_reg0.q\[8\] _06320_ VPWR VGND sg13g2_nor2_1
X_11501_ _05406_ net1840 fp16_sum_pipe.add_renorm0.mantisa\[5\] VPWR VGND sg13g2_nand2_1
X_14220_ _00021_ VGND VPWR _00771_ sipo.shift_reg\[1\] clknet_leaf_21_clk sg13g2_dfrbpq_1
X_11432_ _05364_ VPWR _01056_ VGND net1938 _05363_ sg13g2_o21ai_1
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_11_177 VPWR VGND sg13g2_decap_8
XFILLER_118_0 VPWR VGND sg13g2_decap_8
X_14151_ VPWR _00702_ net131 VGND sg13g2_inv_1
XFILLER_4_811 VPWR VGND sg13g2_decap_8
X_13102_ _06860_ _06791_ _06801_ _06861_ VPWR VGND sg13g2_nand3_1
X_11363_ _05315_ net1812 _05192_ acc_sum.exp_mant_logic0.b\[4\] _05181_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_3_310 VPWR VGND sg13g2_decap_8
X_14082_ VPWR _00633_ net138 VGND sg13g2_inv_1
XFILLER_98_66 VPWR VGND sg13g2_fill_2
X_11294_ acc_sum.reg1en.q\[0\] _05253_ _05046_ _05254_ VPWR VGND sg13g2_nand3_1
XFILLER_65_1010 VPWR VGND sg13g2_decap_4
X_10314_ _04374_ VPWR _01184_ VGND net1919 _04022_ sg13g2_o21ai_1
XFILLER_121_720 VPWR VGND sg13g2_fill_1
XFILLER_79_634 VPWR VGND sg13g2_fill_2
XFILLER_79_612 VPWR VGND sg13g2_decap_8
XFILLER_78_111 VPWR VGND sg13g2_decap_4
X_13033_ _06795_ _06800_ _06801_ VPWR VGND sg13g2_nor2_2
XFILLER_4_888 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
X_10245_ _04315_ _04316_ _04312_ _04317_ VPWR VGND sg13g2_nand3_1
X_10176_ _03611_ _04227_ _04255_ VPWR VGND sg13g2_nor2_1
XFILLER_120_252 VPWR VGND sg13g2_decap_8
XFILLER_93_103 VPWR VGND sg13g2_fill_2
XFILLER_78_177 VPWR VGND sg13g2_decap_8
XFILLER_120_296 VPWR VGND sg13g2_fill_2
XFILLER_66_328 VPWR VGND sg13g2_decap_8
XFILLER_59_380 VPWR VGND sg13g2_fill_2
XFILLER_19_255 VPWR VGND sg13g2_decap_8
X_13935_ VPWR _00486_ net12 VGND sg13g2_inv_1
XFILLER_90_832 VPWR VGND sg13g2_decap_8
XFILLER_47_575 VPWR VGND sg13g2_fill_1
XFILLER_34_225 VPWR VGND sg13g2_decap_4
XFILLER_34_214 VPWR VGND sg13g2_fill_2
X_13866_ VPWR _00417_ net51 VGND sg13g2_inv_1
XFILLER_90_854 VPWR VGND sg13g2_fill_1
X_12817_ _06600_ _06599_ net1959 VPWR VGND sg13g2_nand2_1
XFILLER_34_247 VPWR VGND sg13g2_decap_4
XFILLER_34_236 VPWR VGND sg13g2_decap_8
X_13797_ VPWR _00348_ net81 VGND sg13g2_inv_1
XFILLER_72_1003 VPWR VGND sg13g2_decap_8
XFILLER_50_729 VPWR VGND sg13g2_decap_8
XFILLER_16_973 VPWR VGND sg13g2_decap_8
XFILLER_31_921 VPWR VGND sg13g2_decap_8
X_12748_ fpmul.reg_b_out\[9\] fp16_res_pipe.x2\[9\] net1952 _00919_ VPWR VGND sg13g2_mux2_1
X_12679_ _06490_ _06491_ _06466_ _06492_ VPWR VGND sg13g2_nand3_1
XFILLER_33_1009 VPWR VGND sg13g2_decap_4
XFILLER_8_42 VPWR VGND sg13g2_decap_8
XFILLER_30_453 VPWR VGND sg13g2_fill_1
X_14418_ _00219_ VGND VPWR _00957_ fpmul.reg_a_out\[15\] clknet_leaf_126_clk sg13g2_dfrbpq_1
XFILLER_31_998 VPWR VGND sg13g2_decap_8
X_14349_ _00150_ VGND VPWR _00891_ fpmul.reg_p_out\[13\] clknet_leaf_94_clk sg13g2_dfrbpq_1
XFILLER_7_671 VPWR VGND sg13g2_decap_8
XFILLER_104_709 VPWR VGND sg13g2_fill_2
X_08910_ _03097_ _03096_ VPWR VGND sg13g2_inv_2
XFILLER_112_720 VPWR VGND sg13g2_decap_4
XFILLER_98_932 VPWR VGND sg13g2_decap_8
X_09890_ VPWR _03987_ fp16_res_pipe.seg_reg0.q\[29\] VGND sg13g2_inv_1
XFILLER_33_0 VPWR VGND sg13g2_decap_8
XFILLER_112_775 VPWR VGND sg13g2_decap_8
XFILLER_100_937 VPWR VGND sg13g2_decap_8
XFILLER_84_136 VPWR VGND sg13g2_fill_2
X_08772_ VPWR _02961_ acc_sum.exp_mant_logic0.a\[1\] VGND sg13g2_inv_1
X_07723_ _02030_ net1780 acc_sub.op_sign_logic0.mantisa_a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_66_862 VPWR VGND sg13g2_fill_2
XFILLER_66_851 VPWR VGND sg13g2_decap_8
XFILLER_38_553 VPWR VGND sg13g2_fill_1
X_07654_ _01428_ _01964_ _01965_ VPWR VGND sg13g2_nand2_1
XFILLER_93_681 VPWR VGND sg13g2_fill_2
XFILLER_93_670 VPWR VGND sg13g2_fill_2
XFILLER_81_821 VPWR VGND sg13g2_decap_4
XFILLER_65_372 VPWR VGND sg13g2_fill_2
XFILLER_25_203 VPWR VGND sg13g2_fill_2
XFILLER_25_236 VPWR VGND sg13g2_fill_1
X_07585_ _01898_ VPWR _01899_ VGND _01875_ net1687 sg13g2_o21ai_1
XFILLER_80_375 VPWR VGND sg13g2_decap_8
XFILLER_53_589 VPWR VGND sg13g2_decap_8
XFILLER_43_28 VPWR VGND sg13g2_decap_8
X_09324_ _03477_ _03476_ _03376_ VPWR VGND sg13g2_nand2_1
XFILLER_22_954 VPWR VGND sg13g2_decap_8
X_09255_ VPWR _03409_ fp16_res_pipe.op_sign_logic0.mantisa_b\[0\] VGND sg13g2_inv_1
X_08206_ _02210_ _02227_ _02205_ _02462_ VPWR VGND _02216_ sg13g2_nand4_1
XFILLER_119_363 VPWR VGND sg13g2_fill_2
XFILLER_119_352 VPWR VGND sg13g2_decap_8
X_09186_ _03347_ acc_sum.exp_mant_logic0.b\[5\] VPWR VGND sg13g2_inv_2
XFILLER_111_7 VPWR VGND sg13g2_decap_8
X_08137_ _02272_ _02396_ _02398_ VPWR VGND sg13g2_nor2_1
XFILLER_108_21 VPWR VGND sg13g2_decap_8
X_08068_ VPWR _02334_ _02332_ VGND sg13g2_inv_1
XFILLER_122_528 VPWR VGND sg13g2_fill_2
XFILLER_122_517 VPWR VGND sg13g2_fill_1
Xplace1871 net1870 net1871 VPWR VGND sg13g2_buf_2
Xplace1860 fpmul.reg_a_out\[0\] net1860 VPWR VGND sg13g2_buf_2
XFILLER_1_836 VPWR VGND sg13g2_decap_8
XFILLER_89_965 VPWR VGND sg13g2_decap_8
Xplace1893 acc_sub.reg1en.d\[0\] net1893 VPWR VGND sg13g2_buf_2
Xplace1882 net1881 net1882 VPWR VGND sg13g2_buf_1
XFILLER_0_313 VPWR VGND sg13g2_decap_8
X_10030_ VGND VPWR _04038_ _04051_ _04118_ _04117_ sg13g2_a21oi_1
XFILLER_103_775 VPWR VGND sg13g2_fill_2
XFILLER_0_379 VPWR VGND sg13g2_decap_8
XFILLER_124_42 VPWR VGND sg13g2_decap_8
XFILLER_29_520 VPWR VGND sg13g2_fill_1
XFILLER_29_531 VPWR VGND sg13g2_decap_8
XFILLER_75_158 VPWR VGND sg13g2_fill_2
XFILLER_57_862 VPWR VGND sg13g2_decap_4
XFILLER_56_350 VPWR VGND sg13g2_decap_4
X_11981_ _05835_ _05832_ _05834_ VPWR VGND sg13g2_xnor2_1
X_13720_ VPWR _00271_ net139 VGND sg13g2_inv_1
X_10932_ _04939_ VPWR _01131_ VGND fp16_res_pipe.reg3en.q\[0\] _04929_ sg13g2_o21ai_1
XFILLER_72_854 VPWR VGND sg13g2_fill_2
XFILLER_72_843 VPWR VGND sg13g2_fill_1
XFILLER_71_342 VPWR VGND sg13g2_decap_8
XFILLER_44_556 VPWR VGND sg13g2_fill_1
XFILLER_16_236 VPWR VGND sg13g2_decap_8
XFILLER_16_247 VPWR VGND sg13g2_fill_2
XFILLER_72_898 VPWR VGND sg13g2_fill_1
X_13651_ VPWR _00202_ net110 VGND sg13g2_inv_1
XFILLER_44_567 VPWR VGND sg13g2_decap_8
X_10863_ _04862_ _04874_ _04875_ VPWR VGND sg13g2_nor2_1
XFILLER_31_217 VPWR VGND sg13g2_decap_8
X_13582_ VPWR _00133_ net118 VGND sg13g2_inv_1
X_12602_ _06418_ _06403_ _06405_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_420 VPWR VGND sg13g2_decap_8
XFILLER_13_954 VPWR VGND sg13g2_decap_8
X_10794_ VPWR _04806_ _04805_ VGND sg13g2_inv_1
X_12533_ _06352_ VPWR _00943_ VGND net1954 _05881_ sg13g2_o21ai_1
XFILLER_40_740 VPWR VGND sg13g2_decap_8
XFILLER_9_969 VPWR VGND sg13g2_decap_8
X_14203_ VPWR _00754_ net103 VGND sg13g2_inv_1
X_12464_ _06306_ _06250_ _06152_ VPWR VGND sg13g2_nand2b_1
XFILLER_126_834 VPWR VGND sg13g2_decap_8
XFILLER_125_322 VPWR VGND sg13g2_decap_8
X_11415_ _05354_ net1707 fpdiv.div_out\[1\] VPWR VGND sg13g2_nand2_1
X_12395_ _06223_ _06212_ _06241_ VPWR VGND sg13g2_nor2_1
X_14134_ VPWR _00685_ net89 VGND sg13g2_inv_1
X_11346_ _05299_ net1697 acc_sum.exp_mant_logic0.b\[0\] VPWR VGND sg13g2_nand2_1
X_14065_ VPWR _00616_ net94 VGND sg13g2_inv_1
XFILLER_3_140 VPWR VGND sg13g2_decap_8
XFILLER_98_239 VPWR VGND sg13g2_decap_8
X_13016_ VPWR _06784_ _06783_ VGND sg13g2_inv_1
X_11277_ _05239_ _05237_ _05238_ VPWR VGND sg13g2_nand2_1
XFILLER_67_604 VPWR VGND sg13g2_fill_2
X_10228_ _04300_ _04156_ _04301_ VPWR VGND sg13g2_nor2_1
XFILLER_95_946 VPWR VGND sg13g2_decap_8
XFILLER_0_891 VPWR VGND sg13g2_decap_8
X_10159_ _04240_ _04231_ _04239_ VPWR VGND sg13g2_nand2_1
X_14967_ _00768_ VGND VPWR _01487_ acc_sub.add_renorm0.mantisa\[11\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_1
XFILLER_94_467 VPWR VGND sg13g2_decap_4
XFILLER_82_618 VPWR VGND sg13g2_decap_8
XFILLER_94_489 VPWR VGND sg13g2_fill_2
XFILLER_48_895 VPWR VGND sg13g2_decap_8
XFILLER_48_884 VPWR VGND sg13g2_decap_4
X_14898_ _00699_ VGND VPWR _01418_ acc_sub.op_sign_logic0.mantisa_b\[8\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_2
XFILLER_63_854 VPWR VGND sg13g2_fill_2
X_13918_ VPWR _00469_ net8 VGND sg13g2_inv_1
XFILLER_74_90 VPWR VGND sg13g2_fill_2
XFILLER_50_504 VPWR VGND sg13g2_decap_4
X_13849_ VPWR _00400_ net30 VGND sg13g2_inv_1
XFILLER_22_206 VPWR VGND sg13g2_fill_1
X_07370_ _01722_ VPWR _01469_ VGND net1798 _01721_ sg13g2_o21ai_1
XFILLER_22_239 VPWR VGND sg13g2_decap_8
X_09040_ _03224_ _03225_ _03226_ VPWR VGND sg13g2_nor2b_1
XFILLER_30_283 VPWR VGND sg13g2_fill_2
XFILLER_117_823 VPWR VGND sg13g2_decap_8
XFILLER_116_366 VPWR VGND sg13g2_decap_8
X_09942_ VGND VPWR _04036_ _04024_ _04038_ _04037_ sg13g2_a21oi_1
X_09873_ VGND VPWR _03978_ net1803 _03979_ _03743_ sg13g2_a21oi_1
XFILLER_86_924 VPWR VGND sg13g2_decap_8
X_08824_ _02979_ _02995_ _03011_ VPWR VGND sg13g2_nor2_1
XFILLER_100_723 VPWR VGND sg13g2_decap_8
XFILLER_97_272 VPWR VGND sg13g2_decap_8
XFILLER_57_103 VPWR VGND sg13g2_decap_4
XFILLER_38_28 VPWR VGND sg13g2_decap_8
XFILLER_85_456 VPWR VGND sg13g2_fill_2
X_08755_ _02950_ acc\[7\] net1896 VPWR VGND sg13g2_nand2_1
XFILLER_39_840 VPWR VGND sg13g2_decap_8
X_07706_ _01424_ _02012_ _02013_ VPWR VGND sg13g2_nand2_1
XFILLER_72_117 VPWR VGND sg13g2_decap_8
XFILLER_54_810 VPWR VGND sg13g2_decap_4
XFILLER_38_372 VPWR VGND sg13g2_decap_8
X_08686_ _02757_ _02766_ _02901_ VPWR VGND sg13g2_nor2_1
XFILLER_38_383 VPWR VGND sg13g2_decap_4
XFILLER_54_49 VPWR VGND sg13g2_decap_8
X_07568_ _01882_ _01880_ _01881_ VPWR VGND sg13g2_nand2_1
XFILLER_110_77 VPWR VGND sg13g2_decap_8
X_09307_ _03460_ _03443_ _03459_ VPWR VGND sg13g2_nand2b_1
XFILLER_110_88 VPWR VGND sg13g2_fill_1
XFILLER_108_812 VPWR VGND sg13g2_fill_1
XFILLER_6_906 VPWR VGND sg13g2_decap_8
X_09238_ VPWR _03392_ fp16_res_pipe.op_sign_logic0.mantisa_b\[5\] VGND sg13g2_inv_1
XFILLER_10_968 VPWR VGND sg13g2_decap_8
XFILLER_126_119 VPWR VGND sg13g2_decap_8
XFILLER_119_42 VPWR VGND sg13g2_decap_8
X_09169_ _03336_ acc_sub.x2\[11\] net1904 VPWR VGND sg13g2_nand2_1
XFILLER_119_182 VPWR VGND sg13g2_decap_8
XFILLER_107_355 VPWR VGND sg13g2_fill_1
XFILLER_107_344 VPWR VGND sg13g2_decap_8
X_11200_ _05167_ _05073_ net1661 net1808 _05141_ VPWR VGND sg13g2_a22oi_1
X_12180_ _06025_ _05925_ _06026_ VPWR VGND sg13g2_nor2_1
XFILLER_122_314 VPWR VGND sg13g2_fill_2
X_11131_ _05101_ _05002_ _05100_ VPWR VGND sg13g2_xnor2_1
XFILLER_123_848 VPWR VGND sg13g2_decap_8
XFILLER_122_347 VPWR VGND sg13g2_decap_8
Xplace1690 _03828_ net1690 VPWR VGND sg13g2_buf_2
XFILLER_122_369 VPWR VGND sg13g2_decap_4
XFILLER_95_23 VPWR VGND sg13g2_decap_4
X_11062_ _05009_ _04998_ _05040_ VPWR VGND sg13g2_nor2_1
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_1_677 VPWR VGND sg13g2_fill_1
XFILLER_103_572 VPWR VGND sg13g2_fill_2
XFILLER_95_56 VPWR VGND sg13g2_decap_8
XFILLER_77_935 VPWR VGND sg13g2_fill_2
XFILLER_49_648 VPWR VGND sg13g2_decap_4
X_10013_ _04039_ _04084_ net1689 _04101_ VPWR VGND sg13g2_mux2_1
XFILLER_1_699 VPWR VGND sg13g2_decap_4
X_14821_ _00622_ VGND VPWR _01345_ acc_sum.add_renorm0.mantisa\[10\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_64_607 VPWR VGND sg13g2_fill_1
XFILLER_36_309 VPWR VGND sg13g2_decap_8
XFILLER_63_117 VPWR VGND sg13g2_decap_8
XFILLER_48_169 VPWR VGND sg13g2_fill_2
X_14752_ _00553_ VGND VPWR net1819 acc_sum.reg3en.q\[0\] clknet_leaf_24_clk sg13g2_dfrbpq_2
XFILLER_45_854 VPWR VGND sg13g2_fill_2
X_11964_ _05820_ net1883 fpmul.reg_b_out\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_17_534 VPWR VGND sg13g2_fill_1
XFILLER_72_673 VPWR VGND sg13g2_decap_4
X_11895_ fpmul.seg_reg0.q\[53\] fpmul.reg_a_out\[14\] net1878 _01007_ VPWR VGND sg13g2_mux2_1
X_13703_ VPWR _00254_ net50 VGND sg13g2_inv_1
X_14683_ _00484_ VGND VPWR _01211_ fp16_res_pipe.op_sign_logic0.mantisa_a\[9\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_2
X_10915_ VPWR _04924_ _04874_ VGND sg13g2_inv_1
X_13634_ VPWR _00185_ net59 VGND sg13g2_inv_1
X_10846_ VGND VPWR _04782_ net1825 _04858_ _04857_ sg13g2_a21oi_1
XFILLER_32_537 VPWR VGND sg13g2_decap_8
XFILLER_13_751 VPWR VGND sg13g2_decap_8
X_13565_ VPWR _00116_ net82 VGND sg13g2_inv_1
XFILLER_40_570 VPWR VGND sg13g2_decap_8
XFILLER_8_210 VPWR VGND sg13g2_decap_4
X_10777_ VPWR _04789_ _04788_ VGND sg13g2_inv_1
XFILLER_74_7 VPWR VGND sg13g2_decap_4
X_12516_ VGND VPWR _05367_ net1958 _00951_ _06343_ sg13g2_a21oi_1
X_13496_ VPWR _00047_ net32 VGND sg13g2_inv_1
XFILLER_117_119 VPWR VGND sg13g2_decap_8
X_12447_ _06293_ _05876_ fpmul.seg_reg0.q\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_114_804 VPWR VGND sg13g2_decap_8
XFILLER_5_21 VPWR VGND sg13g2_decap_8
XFILLER_119_1003 VPWR VGND sg13g2_decap_8
XFILLER_113_314 VPWR VGND sg13g2_fill_1
XFILLER_99_515 VPWR VGND sg13g2_decap_4
X_12378_ _06224_ _06212_ _06223_ VPWR VGND sg13g2_nand2_1
XFILLER_5_983 VPWR VGND sg13g2_decap_8
X_14117_ VPWR _00668_ net44 VGND sg13g2_inv_1
XFILLER_125_196 VPWR VGND sg13g2_decap_8
XFILLER_113_325 VPWR VGND sg13g2_fill_2
X_11329_ _05281_ _05282_ _05283_ _05284_ VPWR VGND sg13g2_nor3_1
XFILLER_5_98 VPWR VGND sg13g2_decap_8
XFILLER_68_902 VPWR VGND sg13g2_decap_4
X_14048_ VPWR _00599_ net75 VGND sg13g2_inv_1
XFILLER_79_272 VPWR VGND sg13g2_decap_8
XFILLER_67_434 VPWR VGND sg13g2_decap_8
XFILLER_68_979 VPWR VGND sg13g2_decap_8
XFILLER_67_445 VPWR VGND sg13g2_fill_1
XFILLER_39_158 VPWR VGND sg13g2_fill_2
XFILLER_39_147 VPWR VGND sg13g2_decap_8
XFILLER_54_117 VPWR VGND sg13g2_fill_2
X_08540_ _02764_ _02763_ acc_sum.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_35_331 VPWR VGND sg13g2_decap_8
X_08471_ _02702_ _02672_ _02671_ VPWR VGND sg13g2_xnor2_1
XFILLER_91_982 VPWR VGND sg13g2_decap_8
XFILLER_50_312 VPWR VGND sg13g2_fill_1
X_07353_ VPWR _01711_ acc_sub.add_renorm0.exp\[6\] VGND sg13g2_inv_1
X_07284_ VGND VPWR _01632_ net1665 _01652_ _01651_ sg13g2_a21oi_1
X_09023_ _03209_ _03208_ _03195_ VPWR VGND sg13g2_nand2_1
XFILLER_85_1013 VPWR VGND sg13g2_fill_1
XFILLER_116_152 VPWR VGND sg13g2_decap_8
XFILLER_104_336 VPWR VGND sg13g2_fill_2
XFILLER_49_49 VPWR VGND sg13g2_decap_8
X_09925_ VPWR _04022_ fp16_res_pipe.exp_mant_logic0.b\[9\] VGND sg13g2_inv_1
XFILLER_105_22 VPWR VGND sg13g2_decap_8
XFILLER_98_592 VPWR VGND sg13g2_decap_4
XFILLER_98_570 VPWR VGND sg13g2_decap_4
X_09856_ _03965_ VPWR _01233_ VGND net1820 _03956_ sg13g2_o21ai_1
XFILLER_58_434 VPWR VGND sg13g2_decap_8
X_08807_ _02993_ _02977_ _02994_ VPWR VGND sg13g2_and2_1
XFILLER_59_979 VPWR VGND sg13g2_decap_8
X_09787_ _01238_ _03900_ _03901_ VPWR VGND sg13g2_nand2_1
XFILLER_85_264 VPWR VGND sg13g2_decap_8
XFILLER_74_938 VPWR VGND sg13g2_fill_1
XFILLER_46_618 VPWR VGND sg13g2_decap_4
XFILLER_18_309 VPWR VGND sg13g2_fill_2
X_08738_ _02938_ VPWR _01324_ VGND net1904 _02937_ sg13g2_o21ai_1
XFILLER_27_832 VPWR VGND sg13g2_decap_8
XFILLER_121_21 VPWR VGND sg13g2_decap_8
X_08669_ _02887_ _02743_ _02886_ VPWR VGND sg13g2_xnor2_1
XFILLER_82_982 VPWR VGND sg13g2_decap_8
XFILLER_54_662 VPWR VGND sg13g2_fill_1
XFILLER_26_353 VPWR VGND sg13g2_decap_8
XFILLER_27_876 VPWR VGND sg13g2_decap_8
XFILLER_81_492 VPWR VGND sg13g2_fill_2
XFILLER_81_36 VPWR VGND sg13g2_decap_8
XFILLER_42_857 VPWR VGND sg13g2_decap_4
XFILLER_42_824 VPWR VGND sg13g2_decap_8
X_10700_ _04713_ net1826 fp16_res_pipe.add_renorm0.mantisa\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_121_98 VPWR VGND sg13g2_decap_8
X_10631_ VPWR _04644_ fp16_res_pipe.add_renorm0.mantisa\[7\] VGND sg13g2_inv_1
XFILLER_14_63 VPWR VGND sg13g2_decap_8
XFILLER_127_406 VPWR VGND sg13g2_decap_8
X_13350_ _07049_ net1724 fp16_res_pipe.x2\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_6_703 VPWR VGND sg13g2_fill_1
XFILLER_22_592 VPWR VGND sg13g2_decap_8
X_10562_ VPWR _04593_ fp16_sum_pipe.add_renorm0.exp\[1\] VGND sg13g2_inv_1
XFILLER_108_620 VPWR VGND sg13g2_decap_8
X_13281_ acc\[7\] net1676 _06998_ VPWR VGND sg13g2_nor2_1
X_12301_ _06062_ _06146_ _06147_ VPWR VGND sg13g2_nor2_1
XFILLER_6_725 VPWR VGND sg13g2_fill_1
XFILLER_108_642 VPWR VGND sg13g2_fill_1
X_12232_ _06078_ fpmul.reg_a_out\[6\] net1869 VPWR VGND sg13g2_nand2_1
X_10493_ VPWR _04538_ _04513_ VGND sg13g2_inv_1
XFILLER_108_675 VPWR VGND sg13g2_decap_8
XFILLER_100_0 VPWR VGND sg13g2_decap_4
XFILLER_123_656 VPWR VGND sg13g2_fill_1
XFILLER_123_645 VPWR VGND sg13g2_decap_8
X_12163_ _06009_ _06008_ _05983_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_84 VPWR VGND sg13g2_decap_8
XFILLER_123_689 VPWR VGND sg13g2_fill_1
XFILLER_122_133 VPWR VGND sg13g2_decap_8
X_11114_ VGND VPWR _05083_ _05005_ _05084_ _05004_ sg13g2_a21oi_1
X_12094_ _05940_ _05938_ _05939_ VPWR VGND sg13g2_nand2_1
XFILLER_2_975 VPWR VGND sg13g2_decap_8
XFILLER_77_732 VPWR VGND sg13g2_decap_4
X_11045_ _05024_ _05020_ _05023_ VPWR VGND sg13g2_nand2_2
XFILLER_49_423 VPWR VGND sg13g2_decap_8
XFILLER_49_412 VPWR VGND sg13g2_fill_1
XFILLER_1_485 VPWR VGND sg13g2_decap_8
XFILLER_76_220 VPWR VGND sg13g2_fill_2
XFILLER_65_905 VPWR VGND sg13g2_decap_4
XFILLER_77_787 VPWR VGND sg13g2_decap_8
XFILLER_76_275 VPWR VGND sg13g2_fill_2
XFILLER_76_264 VPWR VGND sg13g2_decap_4
XFILLER_49_489 VPWR VGND sg13g2_decap_8
XFILLER_18_821 VPWR VGND sg13g2_decap_8
X_14804_ _00605_ VGND VPWR _01328_ acc_sum.add_renorm0.exp\[1\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
X_12996_ fpmul.seg_reg0.q\[15\] fpmul.seg_reg0.q\[16\] _06764_ VPWR VGND sg13g2_xor2_1
XFILLER_55_70 VPWR VGND sg13g2_decap_8
X_11947_ _05808_ VPWR _00985_ VGND net1874 _05807_ sg13g2_o21ai_1
X_14735_ _00536_ VGND VPWR _01263_ fp16_res_pipe.add_renorm0.exp\[6\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_1
XFILLER_33_813 VPWR VGND sg13g2_decap_8
XFILLER_17_353 VPWR VGND sg13g2_decap_8
XFILLER_33_846 VPWR VGND sg13g2_decap_8
X_11878_ _05767_ _05766_ VPWR VGND sg13g2_inv_2
XFILLER_60_643 VPWR VGND sg13g2_decap_4
X_14666_ _00467_ VGND VPWR _01194_ fp16_res_pipe.op_sign_logic0.mantisa_b\[3\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_2
XFILLER_32_356 VPWR VGND sg13g2_fill_1
X_13617_ VPWR _00168_ net112 VGND sg13g2_inv_1
X_14597_ _00398_ VGND VPWR _01129_ fp16_res_pipe.y\[8\] clknet_leaf_128_clk sg13g2_dfrbpq_2
XFILLER_20_529 VPWR VGND sg13g2_decap_8
X_10829_ _04841_ fp16_res_pipe.add_renorm0.exp\[0\] _04786_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_367 VPWR VGND sg13g2_decap_8
X_13548_ VPWR _00099_ net88 VGND sg13g2_inv_1
XFILLER_9_530 VPWR VGND sg13g2_fill_1
XFILLER_9_585 VPWR VGND sg13g2_fill_1
X_13479_ VPWR _00030_ net16 VGND sg13g2_inv_1
XFILLER_127_995 VPWR VGND sg13g2_decap_8
XFILLER_126_461 VPWR VGND sg13g2_fill_1
XFILLER_126_450 VPWR VGND sg13g2_decap_8
XFILLER_126_494 VPWR VGND sg13g2_fill_2
XFILLER_113_133 VPWR VGND sg13g2_fill_2
XFILLER_99_367 VPWR VGND sg13g2_fill_1
X_07971_ _02244_ _02241_ _02223_ VPWR VGND sg13g2_nand2_2
X_09710_ VGND VPWR _03795_ _03823_ _03826_ _03825_ sg13g2_a21oi_1
XFILLER_67_220 VPWR VGND sg13g2_decap_8
XFILLER_56_916 VPWR VGND sg13g2_decap_8
X_09641_ VGND VPWR _03711_ _03701_ _03758_ _03706_ sg13g2_a21oi_1
XFILLER_68_798 VPWR VGND sg13g2_decap_4
XFILLER_28_629 VPWR VGND sg13g2_fill_2
X_09572_ _03686_ _03688_ _03685_ _03689_ VPWR VGND sg13g2_nand3_1
XFILLER_83_779 VPWR VGND sg13g2_decap_8
XFILLER_82_256 VPWR VGND sg13g2_fill_2
X_08523_ VPWR _02747_ acc_sum.op_sign_logic0.mantisa_b\[2\] VGND sg13g2_inv_1
XFILLER_70_407 VPWR VGND sg13g2_decap_8
XFILLER_64_982 VPWR VGND sg13g2_decap_8
XFILLER_24_813 VPWR VGND sg13g2_decap_4
XFILLER_82_289 VPWR VGND sg13g2_decap_8
XFILLER_51_621 VPWR VGND sg13g2_decap_8
XFILLER_23_301 VPWR VGND sg13g2_decap_4
XFILLER_23_323 VPWR VGND sg13g2_decap_8
XFILLER_24_824 VPWR VGND sg13g2_decap_8
X_08454_ _02688_ _02652_ fpdiv.divider0.remainder_reg\[12\] VPWR VGND sg13g2_nand2_1
X_07405_ _01745_ acc_sub.exp_mant_logic0.a\[4\] VPWR VGND sg13g2_inv_2
X_08385_ VPWR _02623_ fp16_res_pipe.reg4en.q\[0\] VGND sg13g2_inv_1
XFILLER_52_1012 VPWR VGND sg13g2_fill_2
XFILLER_52_1001 VPWR VGND sg13g2_decap_8
XFILLER_50_175 VPWR VGND sg13g2_fill_1
X_07336_ _01600_ net1744 _01698_ VPWR VGND sg13g2_and2_1
XFILLER_51_28 VPWR VGND sg13g2_decap_8
XFILLER_50_197 VPWR VGND sg13g2_decap_8
XFILLER_109_439 VPWR VGND sg13g2_fill_1
XFILLER_109_428 VPWR VGND sg13g2_decap_8
X_07267_ _01636_ _01584_ _01634_ _01637_ VPWR VGND sg13g2_nand3_1
X_09006_ _03191_ VPWR _03192_ VGND _03149_ _03190_ sg13g2_o21ai_1
X_07198_ _01569_ VPWR _01570_ VGND _01553_ _01567_ sg13g2_o21ai_1
XFILLER_105_601 VPWR VGND sg13g2_fill_1
XFILLER_3_728 VPWR VGND sg13g2_decap_8
XFILLER_3_706 VPWR VGND sg13g2_fill_1
XFILLER_104_111 VPWR VGND sg13g2_fill_2
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_104_155 VPWR VGND sg13g2_decap_8
XFILLER_104_144 VPWR VGND sg13g2_decap_4
XFILLER_120_626 VPWR VGND sg13g2_decap_8
XFILLER_116_54 VPWR VGND sg13g2_decap_8
X_09908_ VPWR _04005_ fp16_res_pipe.exp_mant_logic0.b\[11\] VGND sg13g2_inv_1
X_09839_ _03950_ _03878_ _03840_ VPWR VGND sg13g2_nand2_1
XFILLER_101_873 VPWR VGND sg13g2_decap_8
XFILLER_86_562 VPWR VGND sg13g2_decap_8
XFILLER_47_916 VPWR VGND sg13g2_fill_2
XFILLER_86_595 VPWR VGND sg13g2_decap_8
XFILLER_74_768 VPWR VGND sg13g2_decap_8
XFILLER_74_746 VPWR VGND sg13g2_decap_8
X_12850_ VGND VPWR _04929_ net1911 _06630_ net1924 sg13g2_a21oi_1
X_11801_ _05703_ _05573_ add_result\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_27_662 VPWR VGND sg13g2_fill_1
XFILLER_92_57 VPWR VGND sg13g2_fill_1
X_12781_ _06566_ _06561_ _06565_ VPWR VGND sg13g2_nand2_2
X_14520_ _00321_ VGND VPWR _01056_ fpdiv.reg_a_out\[11\] clknet_leaf_53_clk sg13g2_dfrbpq_1
XFILLER_61_429 VPWR VGND sg13g2_decap_8
XFILLER_15_835 VPWR VGND sg13g2_fill_1
XFILLER_26_161 VPWR VGND sg13g2_fill_1
XFILLER_15_868 VPWR VGND sg13g2_decap_8
X_11732_ _05636_ _04595_ _05583_ VPWR VGND sg13g2_xnor2_1
X_14451_ _00252_ VGND VPWR _00990_ fpmul.seg_reg0.q\[36\] clknet_leaf_122_clk sg13g2_dfrbpq_1
XFILLER_42_676 VPWR VGND sg13g2_decap_8
X_11663_ _05567_ VPWR _05568_ VGND net1836 _05564_ sg13g2_o21ai_1
X_14382_ _00183_ VGND VPWR _00923_ fpmul.reg_b_out\[13\] clknet_leaf_124_clk sg13g2_dfrbpq_2
X_10614_ _04624_ _04626_ _04620_ _04627_ VPWR VGND sg13g2_nand3_1
XFILLER_127_203 VPWR VGND sg13g2_decap_8
XFILLER_10_562 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_130_clk clknet_5_6__leaf_clk clknet_leaf_130_clk VPWR VGND sg13g2_buf_8
X_10545_ _04582_ fp16_sum_pipe.seg_reg0.q\[29\] net1845 VPWR VGND sg13g2_nand2_1
XFILLER_109_984 VPWR VGND sg13g2_decap_8
X_13264_ acc\[11\] net1679 _06985_ VPWR VGND sg13g2_nor2_1
X_10476_ VGND VPWR _04522_ _04391_ _04523_ _04452_ sg13g2_a21oi_1
XFILLER_124_921 VPWR VGND sg13g2_decap_8
XFILLER_123_420 VPWR VGND sg13g2_decap_8
X_12215_ _06061_ _06060_ _05977_ VPWR VGND sg13g2_nand2_1
X_13195_ VPWR _06931_ sipo.shift_reg\[6\] VGND sg13g2_inv_1
XFILLER_123_464 VPWR VGND sg13g2_fill_2
XFILLER_111_604 VPWR VGND sg13g2_fill_1
X_12146_ _05992_ _05991_ _05785_ VPWR VGND sg13g2_nand2_1
XFILLER_124_998 VPWR VGND sg13g2_decap_8
XFILLER_123_486 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_77_551 VPWR VGND sg13g2_decap_8
X_12077_ _05923_ _05922_ _05910_ VPWR VGND sg13g2_nand2_1
XFILLER_49_220 VPWR VGND sg13g2_decap_8
XFILLER_77_562 VPWR VGND sg13g2_fill_2
XFILLER_64_201 VPWR VGND sg13g2_fill_2
X_11028_ acc_sum.exp_mant_logic0.a\[13\] _03331_ _05007_ VPWR VGND sg13g2_nor2_1
XFILLER_37_415 VPWR VGND sg13g2_decap_4
XFILLER_2_77 VPWR VGND sg13g2_decap_8
XFILLER_77_595 VPWR VGND sg13g2_fill_1
XFILLER_49_286 VPWR VGND sg13g2_decap_4
XFILLER_46_971 VPWR VGND sg13g2_decap_8
XFILLER_18_651 VPWR VGND sg13g2_decap_8
X_12979_ fpmul.reg_p_out\[15\] fpmul.result\[15\] net1861 _00893_ VPWR VGND sg13g2_mux2_1
XFILLER_52_429 VPWR VGND sg13g2_fill_2
XFILLER_17_150 VPWR VGND sg13g2_fill_1
XFILLER_33_621 VPWR VGND sg13g2_decap_8
XFILLER_17_183 VPWR VGND sg13g2_decap_8
X_14718_ _00519_ VGND VPWR _01246_ fp16_res_pipe.exp_mant_logic0.a\[5\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_14649_ _00450_ VGND VPWR _01177_ fp16_res_pipe.exp_mant_logic0.b\[2\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_2
X_08170_ _02429_ _02378_ fp16_sum_pipe.exp_mant_logic0.a\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_32_186 VPWR VGND sg13g2_decap_4
XFILLER_119_737 VPWR VGND sg13g2_decap_8
XFILLER_118_203 VPWR VGND sg13g2_decap_8
X_07121_ _01494_ acc_sub.op_sign_logic0.s_a acc_sub.op_sign_logic0.s_b VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_121_clk clknet_5_11__leaf_clk clknet_leaf_121_clk VPWR VGND sg13g2_buf_8
XFILLER_106_409 VPWR VGND sg13g2_fill_1
XFILLER_63_0 VPWR VGND sg13g2_decap_4
XFILLER_127_792 VPWR VGND sg13g2_decap_8
XFILLER_126_280 VPWR VGND sg13g2_decap_8
XFILLER_115_921 VPWR VGND sg13g2_decap_8
XFILLER_114_431 VPWR VGND sg13g2_decap_8
XFILLER_99_153 VPWR VGND sg13g2_fill_1
XFILLER_115_998 VPWR VGND sg13g2_decap_8
XFILLER_99_186 VPWR VGND sg13g2_fill_2
XFILLER_99_164 VPWR VGND sg13g2_decap_8
XFILLER_87_315 VPWR VGND sg13g2_decap_8
XFILLER_102_648 VPWR VGND sg13g2_fill_2
X_07954_ _02228_ _02227_ fp16_sum_pipe.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
X_07885_ _02169_ VPWR _01401_ VGND net1895 _01813_ sg13g2_o21ai_1
XFILLER_101_158 VPWR VGND sg13g2_decap_4
XFILLER_56_713 VPWR VGND sg13g2_decap_8
XFILLER_29_927 VPWR VGND sg13g2_decap_8
X_09624_ _03740_ VPWR _03741_ VGND _03734_ _03739_ sg13g2_o21ai_1
XFILLER_46_28 VPWR VGND sg13g2_decap_8
X_09555_ VPWR _03672_ _03671_ VGND sg13g2_inv_1
X_08506_ acc_sum.op_sign_logic0.mantisa_a\[9\] acc_sum.op_sign_logic0.mantisa_b\[9\]
+ _02730_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_963 VPWR VGND sg13g2_decap_8
X_09486_ _03608_ VPWR _01246_ VGND net1917 _03607_ sg13g2_o21ai_1
X_08437_ _02670_ VPWR _02671_ VGND fpdiv.divider0.divisor_reg\[7\] _02658_ sg13g2_o21ai_1
XFILLER_51_473 VPWR VGND sg13g2_decap_4
X_08368_ instr\[3\] instr\[2\] _02611_ VPWR VGND sg13g2_nor2_1
X_07319_ net1744 _01604_ _01682_ _01683_ VPWR VGND sg13g2_nand3_1
XFILLER_109_225 VPWR VGND sg13g2_fill_1
X_08299_ _02459_ _02427_ _02546_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_112_clk clknet_5_9__leaf_clk clknet_leaf_112_clk VPWR VGND sg13g2_buf_8
XFILLER_11_42 VPWR VGND sg13g2_decap_8
X_10330_ _04382_ VPWR _01176_ VGND net1915 _04354_ sg13g2_o21ai_1
XFILLER_127_42 VPWR VGND sg13g2_decap_8
XFILLER_124_217 VPWR VGND sg13g2_decap_8
XFILLER_106_943 VPWR VGND sg13g2_decap_8
XFILLER_105_420 VPWR VGND sg13g2_fill_2
XFILLER_3_525 VPWR VGND sg13g2_decap_8
X_10261_ _04328_ _04331_ _04332_ VPWR VGND sg13g2_nor2_1
X_12000_ _05854_ fpmul.reg_a_out\[12\] fpmul.reg_b_out\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_121_924 VPWR VGND sg13g2_decap_8
XFILLER_105_486 VPWR VGND sg13g2_fill_2
XFILLER_87_46 VPWR VGND sg13g2_decap_4
X_10192_ net1831 _04268_ net1689 _04270_ VPWR VGND sg13g2_nand3_1
XFILLER_120_456 VPWR VGND sg13g2_decap_8
XFILLER_120_489 VPWR VGND sg13g2_decap_8
X_13951_ VPWR _00502_ net98 VGND sg13g2_inv_1
XFILLER_101_692 VPWR VGND sg13g2_fill_2
XFILLER_87_893 VPWR VGND sg13g2_decap_8
X_12902_ _06678_ _06677_ net1962 VPWR VGND sg13g2_nand2_1
XFILLER_74_565 VPWR VGND sg13g2_decap_8
XFILLER_46_267 VPWR VGND sg13g2_decap_4
X_13882_ VPWR _00433_ net48 VGND sg13g2_inv_1
X_12833_ _06613_ _06614_ _06604_ _00906_ VPWR VGND sg13g2_nand3_1
X_12764_ VGND VPWR net1923 add_result\[15\] _06549_ net1941 sg13g2_a21oi_1
XFILLER_15_654 VPWR VGND sg13g2_fill_2
XFILLER_99_9 VPWR VGND sg13g2_fill_1
X_14503_ _00304_ VGND VPWR _01039_ fpdiv.reg_b_out\[10\] clknet_leaf_91_clk sg13g2_dfrbpq_2
XFILLER_43_985 VPWR VGND sg13g2_fill_1
X_11715_ _05617_ _05618_ _05619_ VPWR VGND sg13g2_nor2_1
X_12695_ VPWR _06504_ _06432_ VGND sg13g2_inv_1
XFILLER_14_197 VPWR VGND sg13g2_decap_8
X_14434_ _00235_ VGND VPWR _00973_ fpmul.seg_reg0.q\[19\] clknet_leaf_96_clk sg13g2_dfrbpq_1
X_11646_ _05551_ _05550_ VPWR VGND sg13g2_inv_2
XFILLER_30_668 VPWR VGND sg13g2_decap_4
X_14365_ _00166_ VGND VPWR _00907_ _00018_ clknet_leaf_87_clk sg13g2_dfrbpq_1
Xclkbuf_leaf_103_clk clknet_5_14__leaf_clk clknet_leaf_103_clk VPWR VGND sg13g2_buf_8
XFILLER_11_882 VPWR VGND sg13g2_decap_8
X_11577_ VPWR _05482_ _05477_ VGND sg13g2_inv_1
X_14296_ _00097_ VGND VPWR _00840_ acc\[6\] clknet_leaf_45_clk sg13g2_dfrbpq_2
X_13316_ acc\[0\] _07025_ net1678 _00834_ VPWR VGND sg13g2_mux2_1
XFILLER_7_853 VPWR VGND sg13g2_decap_8
XFILLER_6_330 VPWR VGND sg13g2_decap_8
X_10528_ VGND VPWR _04567_ net1849 _01164_ _04568_ sg13g2_a21oi_1
XFILLER_115_217 VPWR VGND sg13g2_decap_8
X_13247_ _06971_ _02578_ acc_sub.y\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_108_291 VPWR VGND sg13g2_decap_8
X_10459_ VGND VPWR _04506_ _04423_ _04507_ _04422_ sg13g2_a21oi_1
XFILLER_124_795 VPWR VGND sg13g2_decap_8
X_13178_ _06919_ VPWR _00866_ VGND _06918_ net1715 sg13g2_o21ai_1
XFILLER_123_294 VPWR VGND sg13g2_decap_8
XFILLER_112_957 VPWR VGND sg13g2_decap_8
X_12129_ _05966_ _05970_ _05975_ VPWR VGND sg13g2_nor2_1
XFILLER_97_679 VPWR VGND sg13g2_fill_2
XFILLER_42_1011 VPWR VGND sg13g2_fill_2
XFILLER_77_370 VPWR VGND sg13g2_fill_2
XFILLER_65_521 VPWR VGND sg13g2_fill_2
XFILLER_38_724 VPWR VGND sg13g2_fill_2
X_07670_ _01747_ _01979_ _01980_ VPWR VGND sg13g2_nor2_1
XFILLER_26_919 VPWR VGND sg13g2_decap_8
XFILLER_65_576 VPWR VGND sg13g2_decap_4
XFILLER_18_470 VPWR VGND sg13g2_decap_8
XFILLER_19_971 VPWR VGND sg13g2_decap_8
X_09340_ VGND VPWR _03491_ _03425_ _03492_ _03422_ sg13g2_a21oi_1
XFILLER_34_996 VPWR VGND sg13g2_decap_8
X_09271_ _03422_ _03424_ _03425_ VPWR VGND sg13g2_nor2_2
XFILLER_21_602 VPWR VGND sg13g2_decap_8
XFILLER_33_440 VPWR VGND sg13g2_decap_4
XFILLER_33_462 VPWR VGND sg13g2_decap_4
X_08222_ _02477_ net1638 _02474_ VPWR VGND sg13g2_nand2b_1
XFILLER_119_523 VPWR VGND sg13g2_decap_8
X_08153_ _02413_ fp16_sum_pipe.exp_mant_logic0.a\[4\] net1658 net1691 fp16_sum_pipe.exp_mant_logic0.a\[0\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_119_567 VPWR VGND sg13g2_fill_1
XFILLER_9_190 VPWR VGND sg13g2_decap_4
X_08084_ _02345_ _02349_ _02340_ _02350_ VPWR VGND sg13g2_nand3_1
XFILLER_115_795 VPWR VGND sg13g2_decap_8
X_08986_ acc_sub.add_renorm0.exp\[2\] _03146_ _03172_ VPWR VGND sg13g2_nor2_1
XFILLER_103_946 VPWR VGND sg13g2_decap_8
XFILLER_88_657 VPWR VGND sg13g2_decap_8
XFILLER_87_112 VPWR VGND sg13g2_decap_8
XFILLER_102_456 VPWR VGND sg13g2_fill_1
XFILLER_87_167 VPWR VGND sg13g2_decap_8
XFILLER_69_871 VPWR VGND sg13g2_fill_1
X_07937_ _02209_ _02211_ _02212_ VPWR VGND sg13g2_nor2_1
XFILLER_75_329 VPWR VGND sg13g2_decap_8
XFILLER_68_381 VPWR VGND sg13g2_decap_8
XFILLER_56_521 VPWR VGND sg13g2_decap_4
XFILLER_29_735 VPWR VGND sg13g2_decap_8
X_07868_ _02161_ net1885 acc_sub.x2\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_83_340 VPWR VGND sg13g2_fill_2
XFILLER_17_919 VPWR VGND sg13g2_decap_8
XFILLER_113_77 VPWR VGND sg13g2_decap_8
X_09607_ _03724_ net1806 acc_sum.add_renorm0.mantisa\[10\] VPWR VGND sg13g2_nand2_1
X_07799_ _02095_ _02097_ _02098_ VPWR VGND sg13g2_nor2_1
XFILLER_83_384 VPWR VGND sg13g2_fill_2
XFILLER_73_15 VPWR VGND sg13g2_decap_8
X_09538_ _03655_ acc_sum.add_renorm0.mantisa\[4\] _03621_ VPWR VGND sg13g2_xnor2_1
XFILLER_71_535 VPWR VGND sg13g2_fill_1
XFILLER_25_952 VPWR VGND sg13g2_decap_8
XFILLER_12_613 VPWR VGND sg13g2_decap_4
XFILLER_19_1013 VPWR VGND sg13g2_fill_1
XFILLER_52_793 VPWR VGND sg13g2_fill_2
X_09469_ VPWR _03597_ fp16_res_pipe.exp_mant_logic0.a\[10\] VGND sg13g2_inv_1
XFILLER_11_112 VPWR VGND sg13g2_fill_1
X_11500_ VPWR _05405_ _05404_ VGND sg13g2_inv_1
XFILLER_24_484 VPWR VGND sg13g2_decap_8
X_12480_ _06319_ _06151_ _06250_ VPWR VGND sg13g2_xnor2_1
XFILLER_51_292 VPWR VGND sg13g2_decap_8
XFILLER_40_966 VPWR VGND sg13g2_decap_8
XFILLER_8_628 VPWR VGND sg13g2_fill_2
XFILLER_7_105 VPWR VGND sg13g2_decap_8
X_11431_ _05364_ acc_sub.x2\[11\] net1938 VPWR VGND sg13g2_nand2_1
XFILLER_40_999 VPWR VGND sg13g2_decap_8
X_14150_ VPWR _00701_ net132 VGND sg13g2_inv_1
X_11362_ _05314_ _05227_ _05253_ net1811 _05211_ VPWR VGND sg13g2_a22oi_1
XFILLER_22_63 VPWR VGND sg13g2_decap_8
X_13101_ _06771_ VPWR _06860_ VGND _06774_ _06788_ sg13g2_o21ai_1
X_10313_ _04374_ net1920 fp16_res_pipe.x2\[9\] VPWR VGND sg13g2_nand2_1
X_14081_ VPWR _00632_ net138 VGND sg13g2_inv_1
XFILLER_106_751 VPWR VGND sg13g2_decap_8
XFILLER_98_45 VPWR VGND sg13g2_decap_8
X_11293_ _05252_ _05253_ VPWR VGND sg13g2_inv_4
XFILLER_4_867 VPWR VGND sg13g2_decap_8
X_13032_ _06799_ _06777_ _06800_ VPWR VGND sg13g2_and2_1
X_10244_ _04316_ net1830 _04177_ fp16_res_pipe.exp_mant_logic0.b\[3\] net1643 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_120_231 VPWR VGND sg13g2_decap_8
XFILLER_3_399 VPWR VGND sg13g2_decap_8
X_10175_ _01203_ _04253_ _04254_ VPWR VGND sg13g2_nand2_1
XFILLER_94_605 VPWR VGND sg13g2_fill_2
XFILLER_121_798 VPWR VGND sg13g2_decap_8
XFILLER_93_126 VPWR VGND sg13g2_fill_1
XFILLER_75_874 VPWR VGND sg13g2_decap_8
XFILLER_47_82 VPWR VGND sg13g2_decap_8
X_13934_ VPWR _00485_ net11 VGND sg13g2_inv_1
XFILLER_19_234 VPWR VGND sg13g2_decap_8
XFILLER_90_811 VPWR VGND sg13g2_decap_8
XFILLER_75_896 VPWR VGND sg13g2_decap_8
X_13865_ VPWR _00416_ net56 VGND sg13g2_inv_1
XFILLER_34_204 VPWR VGND sg13g2_fill_1
X_12816_ VPWR _06599_ fpmul.reg_p_out\[13\] VGND sg13g2_inv_1
XFILLER_62_557 VPWR VGND sg13g2_decap_8
XFILLER_35_749 VPWR VGND sg13g2_decap_8
XFILLER_16_952 VPWR VGND sg13g2_decap_8
XFILLER_63_70 VPWR VGND sg13g2_fill_2
X_13796_ VPWR _00347_ net20 VGND sg13g2_inv_1
XFILLER_43_771 VPWR VGND sg13g2_fill_2
XFILLER_31_900 VPWR VGND sg13g2_decap_8
XFILLER_63_81 VPWR VGND sg13g2_decap_8
X_12747_ fpmul.reg_b_out\[10\] fp16_res_pipe.x2\[10\] net1952 _00920_ VPWR VGND sg13g2_mux2_1
XFILLER_43_793 VPWR VGND sg13g2_decap_8
XFILLER_15_484 VPWR VGND sg13g2_decap_8
X_12678_ _06491_ _06464_ _06417_ VPWR VGND sg13g2_nand2_1
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_31_977 VPWR VGND sg13g2_decap_8
X_14417_ _00218_ VGND VPWR _00956_ fpmul.reg_a_out\[14\] clknet_leaf_125_clk sg13g2_dfrbpq_2
X_11629_ _05534_ _05532_ _05521_ VPWR VGND sg13g2_nand2_1
XFILLER_8_98 VPWR VGND sg13g2_decap_8
X_14348_ _00149_ VGND VPWR _00890_ fpmul.reg_p_out\[12\] clknet_leaf_94_clk sg13g2_dfrbpq_1
X_14279_ _00080_ VGND VPWR _00830_ fp16_res_pipe.x2\[12\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_6_182 VPWR VGND sg13g2_decap_8
XFILLER_124_570 VPWR VGND sg13g2_decap_8
X_08840_ _03026_ VPWR _03027_ VGND _03024_ acc_sub.add_renorm0.mantisa\[4\] sg13g2_o21ai_1
XFILLER_112_754 VPWR VGND sg13g2_decap_8
XFILLER_100_916 VPWR VGND sg13g2_decap_8
XFILLER_98_988 VPWR VGND sg13g2_decap_8
XFILLER_85_616 VPWR VGND sg13g2_decap_8
XFILLER_69_156 VPWR VGND sg13g2_decap_4
XFILLER_26_0 VPWR VGND sg13g2_decap_8
XFILLER_84_115 VPWR VGND sg13g2_decap_8
X_08771_ _02960_ VPWR _01313_ VGND net1899 _02959_ sg13g2_o21ai_1
X_07722_ _02029_ _02028_ _01944_ VPWR VGND sg13g2_nand2_1
XFILLER_81_800 VPWR VGND sg13g2_decap_8
X_07653_ _01965_ acc_sub.exp_mant_logic0.a\[4\] net1672 acc_sub.op_sign_logic0.mantisa_a\[7\]
+ net1780 VPWR VGND sg13g2_a22oi_1
XFILLER_65_362 VPWR VGND sg13g2_fill_1
XFILLER_53_502 VPWR VGND sg13g2_fill_2
XFILLER_38_587 VPWR VGND sg13g2_decap_8
XFILLER_26_716 VPWR VGND sg13g2_decap_4
X_07584_ _01898_ net1687 _01889_ VPWR VGND sg13g2_nand2_1
XFILLER_53_568 VPWR VGND sg13g2_decap_8
X_09323_ _03475_ VPWR _03476_ VGND _03370_ _03434_ sg13g2_o21ai_1
XFILLER_80_398 VPWR VGND sg13g2_decap_8
XFILLER_21_421 VPWR VGND sg13g2_decap_8
XFILLER_22_933 VPWR VGND sg13g2_decap_8
X_09254_ _03408_ _03402_ _03407_ VPWR VGND sg13g2_nand2_1
X_09185_ _03346_ VPWR _01285_ VGND net1905 _03345_ sg13g2_o21ai_1
X_08205_ _02459_ _02460_ _02458_ _02461_ VPWR VGND sg13g2_nand3_1
XFILLER_4_119 VPWR VGND sg13g2_decap_8
Xplace1872 net1871 net1872 VPWR VGND sg13g2_buf_2
Xplace1861 fpmul.reg2en.q\[0\] net1861 VPWR VGND sg13g2_buf_2
Xplace1850 fp16_sum_pipe.reg3en.q\[0\] net1850 VPWR VGND sg13g2_buf_2
XFILLER_1_815 VPWR VGND sg13g2_decap_8
XFILLER_108_88 VPWR VGND sg13g2_decap_4
Xplace1894 net1893 net1894 VPWR VGND sg13g2_buf_1
XFILLER_89_944 VPWR VGND sg13g2_decap_8
Xplace1883 net1882 net1883 VPWR VGND sg13g2_buf_2
XFILLER_124_21 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_decap_8
XFILLER_0_358 VPWR VGND sg13g2_decap_8
X_08969_ VPWR _03155_ _03154_ VGND sg13g2_inv_1
XFILLER_102_286 VPWR VGND sg13g2_fill_2
XFILLER_124_98 VPWR VGND sg13g2_decap_8
X_11980_ fpmul.reg_b_out\[10\] fpmul.reg_a_out\[10\] _05834_ VPWR VGND sg13g2_xor2_1
XFILLER_57_896 VPWR VGND sg13g2_decap_8
X_10931_ _04897_ _04938_ _04936_ _04939_ VPWR VGND sg13g2_nand3_1
XFILLER_84_693 VPWR VGND sg13g2_decap_8
XFILLER_17_63 VPWR VGND sg13g2_decap_8
X_13650_ VPWR _00201_ net110 VGND sg13g2_inv_1
XFILLER_16_259 VPWR VGND sg13g2_decap_8
XFILLER_25_760 VPWR VGND sg13g2_decap_8
X_10862_ _04874_ _04871_ _04873_ VPWR VGND sg13g2_nand2_1
XFILLER_32_708 VPWR VGND sg13g2_fill_1
X_13581_ VPWR _00132_ net114 VGND sg13g2_inv_1
X_12601_ _06417_ _06406_ _06396_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_410 VPWR VGND sg13g2_fill_2
XFILLER_13_933 VPWR VGND sg13g2_decap_8
X_10793_ _04804_ _04777_ _04805_ VPWR VGND sg13g2_and2_1
XFILLER_25_793 VPWR VGND sg13g2_decap_8
X_12532_ _06352_ acc_sub.x2\[1\] net1955 VPWR VGND sg13g2_nand2_1
X_12463_ _06305_ _06020_ _06061_ VPWR VGND sg13g2_nand2_1
XFILLER_40_785 VPWR VGND sg13g2_decap_8
XFILLER_8_425 VPWR VGND sg13g2_decap_8
XFILLER_9_948 VPWR VGND sg13g2_decap_8
XFILLER_12_476 VPWR VGND sg13g2_decap_8
XFILLER_33_84 VPWR VGND sg13g2_fill_2
XFILLER_126_813 VPWR VGND sg13g2_decap_8
X_14202_ VPWR _00753_ net104 VGND sg13g2_inv_1
X_11414_ VPWR _05353_ fpdiv.div_out\[0\] VGND sg13g2_inv_1
XFILLER_8_469 VPWR VGND sg13g2_decap_8
XFILLER_125_301 VPWR VGND sg13g2_decap_8
X_12394_ VGND VPWR _06234_ _06238_ _06240_ _06239_ sg13g2_a21oi_1
XFILLER_99_708 VPWR VGND sg13g2_decap_8
X_14133_ VPWR _00684_ net102 VGND sg13g2_inv_1
X_11345_ _05298_ net1656 acc_sum.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_98_218 VPWR VGND sg13g2_decap_8
X_14064_ VPWR _00615_ net94 VGND sg13g2_inv_1
X_11276_ _05238_ net1810 _05192_ acc_sum.exp_mant_logic0.a\[3\] net1653 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_4_664 VPWR VGND sg13g2_decap_8
X_13015_ _06313_ net1853 _06782_ _06783_ VPWR VGND sg13g2_a21o_1
XFILLER_3_196 VPWR VGND sg13g2_decap_8
X_10227_ _04300_ fp16_res_pipe.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_inv_2
XFILLER_95_903 VPWR VGND sg13g2_fill_2
XFILLER_58_92 VPWR VGND sg13g2_decap_8
XFILLER_58_81 VPWR VGND sg13g2_decap_8
XFILLER_0_870 VPWR VGND sg13g2_decap_8
X_10158_ _04236_ _04238_ _04239_ VPWR VGND sg13g2_nor2_1
X_14966_ _00767_ VGND VPWR _01486_ acc_sub.add_renorm0.mantisa\[10\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_2
XFILLER_48_863 VPWR VGND sg13g2_decap_8
X_10089_ _04174_ _04165_ net1827 VPWR VGND sg13g2_nand2_1
XFILLER_75_660 VPWR VGND sg13g2_fill_1
X_13917_ VPWR _00468_ net8 VGND sg13g2_inv_1
X_14897_ _00698_ VGND VPWR _01417_ acc_sub.op_sign_logic0.mantisa_b\[7\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_2
XFILLER_63_833 VPWR VGND sg13g2_decap_8
XFILLER_62_332 VPWR VGND sg13g2_decap_8
XFILLER_47_395 VPWR VGND sg13g2_decap_8
XFILLER_62_376 VPWR VGND sg13g2_decap_4
X_13848_ VPWR _00399_ net31 VGND sg13g2_inv_1
X_13779_ VPWR _00330_ net137 VGND sg13g2_inv_1
XFILLER_50_527 VPWR VGND sg13g2_decap_8
XFILLER_16_771 VPWR VGND sg13g2_fill_1
XFILLER_15_281 VPWR VGND sg13g2_decap_8
XFILLER_30_251 VPWR VGND sg13g2_decap_4
XFILLER_31_774 VPWR VGND sg13g2_decap_8
XFILLER_31_785 VPWR VGND sg13g2_fill_2
XFILLER_117_802 VPWR VGND sg13g2_decap_8
Xclkbuf_4_4_0_clk clknet_0_clk clknet_4_4_0_clk VPWR VGND sg13g2_buf_8
XFILLER_117_879 VPWR VGND sg13g2_decap_8
XFILLER_116_323 VPWR VGND sg13g2_fill_2
XFILLER_7_491 VPWR VGND sg13g2_decap_8
XFILLER_89_207 VPWR VGND sg13g2_fill_1
X_09941_ VPWR _04037_ _04023_ VGND sg13g2_inv_1
XFILLER_112_551 VPWR VGND sg13g2_fill_2
X_09872_ _03975_ _03976_ _03974_ _03978_ VPWR VGND _03977_ sg13g2_nand4_1
XFILLER_98_752 VPWR VGND sg13g2_decap_8
XFILLER_86_903 VPWR VGND sg13g2_decap_8
X_08823_ _02990_ _03009_ _03010_ VPWR VGND sg13g2_nor2_2
XFILLER_100_713 VPWR VGND sg13g2_decap_4
XFILLER_98_796 VPWR VGND sg13g2_decap_4
XFILLER_100_746 VPWR VGND sg13g2_fill_1
X_08754_ _02949_ acc_sum.exp_mant_logic0.a\[7\] VPWR VGND sg13g2_inv_2
XFILLER_73_608 VPWR VGND sg13g2_fill_1
XFILLER_57_148 VPWR VGND sg13g2_decap_8
X_07705_ _02013_ acc_sub.exp_mant_logic0.a\[0\] net1672 acc_sub.op_sign_logic0.mantisa_a\[3\]
+ net1779 VPWR VGND sg13g2_a22oi_1
XFILLER_39_896 VPWR VGND sg13g2_decap_8
X_08685_ VGND VPWR _02899_ net1817 _01339_ _02900_ sg13g2_a21oi_1
Xclkbuf_leaf_92_clk clknet_5_12__leaf_clk clknet_leaf_92_clk VPWR VGND sg13g2_buf_8
XFILLER_54_844 VPWR VGND sg13g2_fill_1
XFILLER_54_28 VPWR VGND sg13g2_decap_8
X_07636_ _01939_ _01905_ _01949_ VPWR VGND sg13g2_nor2_2
XFILLER_81_674 VPWR VGND sg13g2_fill_1
XFILLER_53_354 VPWR VGND sg13g2_decap_4
XFILLER_14_708 VPWR VGND sg13g2_decap_8
X_07567_ VPWR _01881_ _01815_ VGND sg13g2_inv_1
XFILLER_110_56 VPWR VGND sg13g2_decap_8
X_09306_ _03459_ fp16_res_pipe.op_sign_logic0.mantisa_a\[0\] fp16_res_pipe.op_sign_logic0.mantisa_b\[0\]
+ VPWR VGND sg13g2_nand2_1
X_07498_ _01821_ _01802_ _01820_ VPWR VGND sg13g2_nand2_2
XFILLER_70_49 VPWR VGND sg13g2_fill_1
XFILLER_70_38 VPWR VGND sg13g2_decap_8
X_09237_ VPWR _03391_ _03390_ VGND sg13g2_inv_1
XFILLER_108_802 VPWR VGND sg13g2_fill_1
XFILLER_10_947 VPWR VGND sg13g2_decap_8
XFILLER_119_161 VPWR VGND sg13g2_decap_8
XFILLER_119_21 VPWR VGND sg13g2_decap_8
XFILLER_108_824 VPWR VGND sg13g2_fill_2
XFILLER_107_301 VPWR VGND sg13g2_decap_8
X_09168_ VPWR _03335_ acc_sum.exp_mant_logic0.b\[11\] VGND sg13g2_inv_1
X_09099_ _03281_ VPWR _03282_ VGND net1786 _03279_ sg13g2_o21ai_1
XFILLER_108_857 VPWR VGND sg13g2_decap_8
X_08119_ _02272_ _02380_ _02381_ VPWR VGND sg13g2_nor2_1
XFILLER_123_827 VPWR VGND sg13g2_decap_8
XFILLER_119_98 VPWR VGND sg13g2_decap_8
XFILLER_79_69 VPWR VGND sg13g2_decap_4
X_11130_ _05099_ VPWR _05100_ VGND _05089_ _05046_ sg13g2_o21ai_1
Xplace1680 _05052_ net1680 VPWR VGND sg13g2_buf_2
XFILLER_89_774 VPWR VGND sg13g2_decap_4
X_11061_ _05038_ VPWR _05039_ VGND _05000_ _05037_ sg13g2_o21ai_1
XFILLER_0_133 VPWR VGND sg13g2_decap_8
Xplace1691 _02275_ net1691 VPWR VGND sg13g2_buf_2
XFILLER_88_273 VPWR VGND sg13g2_fill_2
XFILLER_76_413 VPWR VGND sg13g2_fill_1
XFILLER_48_126 VPWR VGND sg13g2_decap_4
X_10012_ _04100_ _03998_ _04099_ VPWR VGND sg13g2_xnor2_1
X_14820_ _00621_ VGND VPWR _01344_ acc_sum.add_renorm0.mantisa\[9\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_77_969 VPWR VGND sg13g2_decap_8
XFILLER_92_939 VPWR VGND sg13g2_decap_8
XFILLER_28_84 VPWR VGND sg13g2_decap_8
X_14751_ _00552_ VGND VPWR acc_sum.reg3en.q\[0\] acc_sum.reg4en.q\[0\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_83_clk clknet_5_26__leaf_clk clknet_leaf_83_clk VPWR VGND sg13g2_buf_8
X_11963_ VPWR _05819_ fpmul.seg_reg0.q\[25\] VGND sg13g2_inv_1
XFILLER_28_95 VPWR VGND sg13g2_fill_2
XFILLER_72_663 VPWR VGND sg13g2_fill_1
XFILLER_60_803 VPWR VGND sg13g2_fill_2
X_11894_ VGND VPWR _05777_ net1876 _01008_ _05778_ sg13g2_a21oi_1
X_13702_ VPWR _00253_ net50 VGND sg13g2_inv_1
X_14682_ _00483_ VGND VPWR _01210_ fp16_res_pipe.op_sign_logic0.mantisa_a\[8\] clknet_leaf_143_clk
+ sg13g2_dfrbpq_2
X_10914_ net1821 _04920_ _04918_ _04923_ VPWR VGND _04922_ sg13g2_nand4_1
XFILLER_60_847 VPWR VGND sg13g2_decap_8
X_13633_ VPWR _00184_ net50 VGND sg13g2_inv_1
X_10845_ net1825 fp16_res_pipe.add_renorm0.exp\[7\] _04857_ VPWR VGND sg13g2_nor2_1
XFILLER_32_527 VPWR VGND sg13g2_fill_2
X_13564_ VPWR _00115_ net82 VGND sg13g2_inv_1
XFILLER_9_712 VPWR VGND sg13g2_decap_8
X_10776_ _04788_ fp16_res_pipe.add_renorm0.exp\[5\] _04779_ VPWR VGND sg13g2_xnor2_1
X_12515_ fpmul.reg_a_out\[9\] net1958 _06343_ VPWR VGND sg13g2_nor2_1
X_13495_ VPWR _00046_ net35 VGND sg13g2_inv_1
XFILLER_12_273 VPWR VGND sg13g2_decap_4
XFILLER_12_295 VPWR VGND sg13g2_decap_8
X_12446_ _06292_ _06291_ net1870 VPWR VGND sg13g2_nand2_1
XFILLER_8_288 VPWR VGND sg13g2_fill_2
X_12377_ _06219_ _06222_ _06223_ VPWR VGND sg13g2_nor2_1
XFILLER_113_304 VPWR VGND sg13g2_fill_1
X_11328_ _03345_ _05148_ _05283_ VPWR VGND sg13g2_nor2_1
XFILLER_5_962 VPWR VGND sg13g2_decap_8
X_14116_ VPWR _00667_ net44 VGND sg13g2_inv_1
XFILLER_125_175 VPWR VGND sg13g2_decap_8
XFILLER_113_348 VPWR VGND sg13g2_fill_2
XFILLER_5_77 VPWR VGND sg13g2_decap_8
XFILLER_4_483 VPWR VGND sg13g2_decap_8
XFILLER_79_251 VPWR VGND sg13g2_decap_8
X_14047_ VPWR _00598_ net76 VGND sg13g2_inv_1
XFILLER_69_80 VPWR VGND sg13g2_fill_2
X_11259_ VPWR _05222_ _05124_ VGND sg13g2_inv_1
XFILLER_122_882 VPWR VGND sg13g2_decap_8
XFILLER_121_370 VPWR VGND sg13g2_decap_8
XFILLER_95_711 VPWR VGND sg13g2_decap_8
XFILLER_68_958 VPWR VGND sg13g2_decap_8
XFILLER_39_126 VPWR VGND sg13g2_decap_8
XFILLER_83_939 VPWR VGND sg13g2_decap_8
X_14949_ _00750_ VGND VPWR _01469_ acc_sub.add_renorm0.exp\[1\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_2
Xclkbuf_leaf_74_clk clknet_5_30__leaf_clk clknet_leaf_74_clk VPWR VGND sg13g2_buf_8
XFILLER_76_991 VPWR VGND sg13g2_decap_8
XFILLER_48_682 VPWR VGND sg13g2_decap_8
XFILLER_35_310 VPWR VGND sg13g2_decap_8
X_08470_ _02701_ VPWR _01355_ VGND net1705 _02700_ sg13g2_o21ai_1
XFILLER_91_961 VPWR VGND sg13g2_decap_8
XFILLER_62_151 VPWR VGND sg13g2_decap_8
XFILLER_39_1005 VPWR VGND sg13g2_decap_8
X_07421_ fpdiv.divider0.state _01755_ _01756_ VPWR VGND sg13g2_nor2_2
XFILLER_62_173 VPWR VGND sg13g2_fill_1
XFILLER_36_899 VPWR VGND sg13g2_decap_8
X_07352_ _01710_ VPWR _01475_ VGND net1797 _01709_ sg13g2_o21ai_1
XFILLER_23_549 VPWR VGND sg13g2_decap_8
X_07283_ _01578_ net1665 _01651_ VPWR VGND sg13g2_nor2_1
X_09022_ VPWR _03208_ _03207_ VGND sg13g2_inv_1
XFILLER_108_109 VPWR VGND sg13g2_decap_4
XFILLER_116_131 VPWR VGND sg13g2_decap_8
XFILLER_117_687 VPWR VGND sg13g2_decap_8
XFILLER_2_409 VPWR VGND sg13g2_decap_8
XFILLER_104_315 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_104_359 VPWR VGND sg13g2_fill_2
XFILLER_104_348 VPWR VGND sg13g2_decap_8
X_09924_ _04021_ _04019_ _04020_ VPWR VGND sg13g2_nand2_1
XFILLER_113_893 VPWR VGND sg13g2_decap_8
X_09855_ _03965_ _03783_ _03964_ VPWR VGND sg13g2_nand2_1
X_08806_ _02993_ _02992_ _01647_ VPWR VGND sg13g2_nand2_1
XFILLER_112_392 VPWR VGND sg13g2_decap_8
XFILLER_85_243 VPWR VGND sg13g2_decap_8
XFILLER_85_232 VPWR VGND sg13g2_fill_1
XFILLER_105_67 VPWR VGND sg13g2_decap_4
X_09786_ _03901_ _03782_ acc_sum.y\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_85_276 VPWR VGND sg13g2_decap_4
XFILLER_27_811 VPWR VGND sg13g2_decap_8
X_08737_ _02938_ acc\[13\] net1901 VPWR VGND sg13g2_nand2_1
X_08668_ VGND VPWR _02884_ _02885_ _02886_ _02831_ sg13g2_a21oi_1
XFILLER_82_961 VPWR VGND sg13g2_decap_8
XFILLER_42_803 VPWR VGND sg13g2_decap_8
XFILLER_26_332 VPWR VGND sg13g2_decap_8
XFILLER_26_343 VPWR VGND sg13g2_decap_8
XFILLER_121_77 VPWR VGND sg13g2_decap_8
X_07619_ _01933_ _01914_ _01918_ VPWR VGND sg13g2_nand2_2
XFILLER_81_471 VPWR VGND sg13g2_decap_8
X_08599_ _02822_ acc_sum.op_sign_logic0.mantisa_a\[2\] acc_sum.op_sign_logic0.mantisa_b\[2\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_14_42 VPWR VGND sg13g2_decap_8
XFILLER_22_582 VPWR VGND sg13g2_fill_1
X_10561_ _04592_ VPWR _01155_ VGND net1844 _04591_ sg13g2_o21ai_1
X_13280_ VPWR VGND acc_sub.y\[7\] _06996_ _02578_ net1742 _06997_ sipo.word\[7\] sg13g2_a221oi_1
X_12300_ VGND VPWR _06135_ _06144_ _06146_ _06145_ sg13g2_a21oi_1
X_10492_ _04536_ net1670 _04537_ VPWR VGND sg13g2_nor2_1
XFILLER_108_654 VPWR VGND sg13g2_decap_8
XFILLER_108_632 VPWR VGND sg13g2_fill_2
X_12231_ _06077_ _06068_ _06076_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_759 VPWR VGND sg13g2_fill_1
XFILLER_5_236 VPWR VGND sg13g2_decap_4
XFILLER_30_63 VPWR VGND sg13g2_decap_8
XFILLER_122_112 VPWR VGND sg13g2_decap_8
XFILLER_107_175 VPWR VGND sg13g2_decap_4
X_12162_ _06008_ _06005_ _06007_ VPWR VGND sg13g2_nand2_1
XFILLER_104_860 VPWR VGND sg13g2_fill_2
X_11113_ VPWR _05083_ _05082_ VGND sg13g2_inv_1
X_12093_ _05932_ _05936_ _05930_ _05939_ VPWR VGND sg13g2_nand3_1
XFILLER_2_954 VPWR VGND sg13g2_decap_8
XFILLER_122_189 VPWR VGND sg13g2_decap_8
XFILLER_104_893 VPWR VGND sg13g2_decap_4
XFILLER_89_593 VPWR VGND sg13g2_decap_8
XFILLER_89_571 VPWR VGND sg13g2_decap_8
X_11044_ _05021_ _05022_ _05023_ VPWR VGND sg13g2_nor2_2
XFILLER_1_464 VPWR VGND sg13g2_decap_8
XFILLER_49_457 VPWR VGND sg13g2_decap_8
XFILLER_65_928 VPWR VGND sg13g2_fill_2
XFILLER_37_608 VPWR VGND sg13g2_decap_4
XFILLER_18_811 VPWR VGND sg13g2_decap_8
XFILLER_92_747 VPWR VGND sg13g2_fill_2
X_14803_ _00604_ VGND VPWR _01327_ acc_sum.add_renorm0.exp\[0\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_2
Xclkbuf_leaf_56_clk clknet_5_28__leaf_clk clknet_leaf_56_clk VPWR VGND sg13g2_buf_8
XFILLER_64_449 VPWR VGND sg13g2_decap_4
X_12995_ VPWR _06763_ _06762_ VGND sg13g2_inv_1
XFILLER_58_991 VPWR VGND sg13g2_fill_1
XFILLER_91_257 VPWR VGND sg13g2_decap_4
XFILLER_91_246 VPWR VGND sg13g2_decap_8
X_11946_ _05808_ net1874 fpmul.reg_b_out\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_44_140 VPWR VGND sg13g2_decap_8
XFILLER_17_332 VPWR VGND sg13g2_decap_4
X_14734_ _00535_ VGND VPWR _01262_ fp16_res_pipe.add_renorm0.exp\[5\] clknet_leaf_131_clk
+ sg13g2_dfrbpq_2
XFILLER_73_983 VPWR VGND sg13g2_decap_4
XFILLER_17_398 VPWR VGND sg13g2_fill_1
XFILLER_18_899 VPWR VGND sg13g2_decap_8
X_11877_ fpdiv.reg1en.q\[0\] fpdiv.divider0.state _05766_ VPWR VGND sg13g2_nor2_1
XFILLER_72_493 VPWR VGND sg13g2_fill_2
X_14665_ _00466_ VGND VPWR _01193_ fp16_res_pipe.op_sign_logic0.mantisa_b\[2\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_1
XFILLER_32_335 VPWR VGND sg13g2_decap_8
X_13616_ VPWR _00167_ net118 VGND sg13g2_inv_1
XFILLER_60_699 VPWR VGND sg13g2_decap_4
X_14596_ _00397_ VGND VPWR _01128_ fp16_res_pipe.y\[7\] clknet_leaf_130_clk sg13g2_dfrbpq_2
X_10828_ _04837_ _04839_ _04840_ VPWR VGND sg13g2_nor2_1
XFILLER_119_919 VPWR VGND sg13g2_decap_8
X_13547_ VPWR _00098_ net88 VGND sg13g2_inv_1
X_10759_ net1835 _04772_ VPWR VGND sg13g2_inv_4
XFILLER_13_593 VPWR VGND sg13g2_decap_8
XFILLER_118_418 VPWR VGND sg13g2_fill_2
X_13478_ VPWR _00029_ net26 VGND sg13g2_inv_1
XFILLER_127_974 VPWR VGND sg13g2_decap_8
X_12429_ _06275_ _06273_ _06274_ VPWR VGND sg13g2_xnor2_1
XFILLER_113_112 VPWR VGND sg13g2_decap_8
XFILLER_5_792 VPWR VGND sg13g2_fill_2
XFILLER_102_808 VPWR VGND sg13g2_fill_2
XFILLER_99_346 VPWR VGND sg13g2_decap_8
XFILLER_87_519 VPWR VGND sg13g2_decap_8
X_07970_ _02243_ VPWR _01390_ VGND net1843 _02226_ sg13g2_o21ai_1
XFILLER_113_167 VPWR VGND sg13g2_decap_4
XFILLER_101_307 VPWR VGND sg13g2_fill_1
XFILLER_95_530 VPWR VGND sg13g2_fill_1
XFILLER_67_210 VPWR VGND sg13g2_fill_2
XFILLER_110_885 VPWR VGND sg13g2_decap_8
X_09640_ _03756_ VPWR _03757_ VGND net1802 _03750_ sg13g2_o21ai_1
X_09571_ _03688_ _03652_ _03687_ _03649_ _03631_ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_47_clk clknet_5_22__leaf_clk clknet_leaf_47_clk VPWR VGND sg13g2_buf_8
X_08522_ VPWR _02746_ _02745_ VGND sg13g2_inv_1
XFILLER_82_268 VPWR VGND sg13g2_fill_2
XFILLER_71_909 VPWR VGND sg13g2_decap_8
X_07404_ _01744_ VPWR _01457_ VGND net1890 _01743_ sg13g2_o21ai_1
XFILLER_51_644 VPWR VGND sg13g2_fill_1
XFILLER_35_195 VPWR VGND sg13g2_fill_2
X_08384_ _02560_ _02619_ _07113_ VPWR VGND sg13g2_nor2_1
XFILLER_50_154 VPWR VGND sg13g2_decap_8
XFILLER_23_368 VPWR VGND sg13g2_decap_4
X_07335_ _01697_ _01564_ _01599_ VPWR VGND sg13g2_nand2b_1
X_07266_ net1783 _01635_ _01636_ VPWR VGND sg13g2_nor2_2
X_09005_ VGND VPWR _03190_ _03149_ _03191_ _03091_ sg13g2_a21oi_1
X_07197_ VGND VPWR _01568_ _01563_ _01569_ _01557_ sg13g2_a21oi_1
XFILLER_118_985 VPWR VGND sg13g2_decap_8
XFILLER_117_495 VPWR VGND sg13g2_decap_4
XFILLER_105_624 VPWR VGND sg13g2_fill_2
XFILLER_2_217 VPWR VGND sg13g2_fill_1
XFILLER_116_33 VPWR VGND sg13g2_decap_8
XFILLER_105_668 VPWR VGND sg13g2_fill_1
XFILLER_99_880 VPWR VGND sg13g2_decap_4
XFILLER_59_711 VPWR VGND sg13g2_fill_2
X_09907_ fp16_res_pipe.exp_mant_logic0.b\[11\] _03595_ _04004_ VPWR VGND sg13g2_nor2_1
XFILLER_98_390 VPWR VGND sg13g2_fill_2
XFILLER_59_755 VPWR VGND sg13g2_decap_8
XFILLER_58_210 VPWR VGND sg13g2_decap_8
XFILLER_47_906 VPWR VGND sg13g2_decap_4
X_09838_ VGND VPWR _03684_ _03851_ _03949_ _03948_ sg13g2_a21oi_1
XFILLER_101_885 VPWR VGND sg13g2_decap_8
XFILLER_74_703 VPWR VGND sg13g2_decap_8
XFILLER_58_276 VPWR VGND sg13g2_decap_8
X_09769_ VGND VPWR _03865_ _03883_ _03885_ _03884_ sg13g2_a21oi_1
Xclkbuf_leaf_38_clk clknet_5_20__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_92_36 VPWR VGND sg13g2_decap_8
XFILLER_92_25 VPWR VGND sg13g2_fill_1
XFILLER_92_14 VPWR VGND sg13g2_decap_8
X_11800_ _05702_ _05699_ _05701_ VPWR VGND sg13g2_nand2_1
X_12780_ net3 _06564_ _06565_ VPWR VGND sg13g2_nor2_1
XFILLER_54_471 VPWR VGND sg13g2_fill_2
XFILLER_54_460 VPWR VGND sg13g2_fill_1
XFILLER_14_313 VPWR VGND sg13g2_decap_8
XFILLER_14_324 VPWR VGND sg13g2_fill_2
XFILLER_25_63 VPWR VGND sg13g2_decap_4
X_11731_ _05635_ _05488_ _05617_ VPWR VGND sg13g2_nand2_1
X_14450_ _00251_ VGND VPWR _00989_ fpmul.seg_reg0.q\[35\] clknet_leaf_122_clk sg13g2_dfrbpq_1
X_11662_ _05566_ _05565_ _05498_ _05567_ VPWR VGND sg13g2_a21o_1
XFILLER_30_806 VPWR VGND sg13g2_decap_8
X_14381_ _00182_ VGND VPWR _00922_ fpmul.reg_b_out\[12\] clknet_leaf_124_clk sg13g2_dfrbpq_2
X_10613_ _04625_ VPWR _04626_ VGND net1826 _04621_ sg13g2_o21ai_1
XFILLER_23_891 VPWR VGND sg13g2_decap_8
X_11593_ _05498_ net1836 VPWR VGND sg13g2_inv_2
X_13332_ VPWR _07037_ sipo.word\[11\] VGND sg13g2_inv_1
X_10544_ _04581_ fp16_sum_pipe.add_renorm0.exp\[7\] VPWR VGND sg13g2_inv_2
XFILLER_41_84 VPWR VGND sg13g2_decap_8
XFILLER_6_523 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_fill_1
XFILLER_10_596 VPWR VGND sg13g2_decap_8
XFILLER_127_259 VPWR VGND sg13g2_decap_8
XFILLER_124_900 VPWR VGND sg13g2_decap_8
XFILLER_109_963 VPWR VGND sg13g2_decap_8
X_13263_ VPWR VGND acc_sum.y\[11\] _06983_ net1729 net1743 _06984_ sipo.word\[11\]
+ sg13g2_a221oi_1
X_10475_ VPWR _04522_ _04450_ VGND sg13g2_inv_1
XFILLER_108_495 VPWR VGND sg13g2_decap_8
XFILLER_108_473 VPWR VGND sg13g2_decap_8
X_12214_ _06060_ _06018_ _06019_ VPWR VGND sg13g2_nand2_1
X_13194_ _06930_ VPWR _00861_ VGND _06929_ net1712 sg13g2_o21ai_1
XFILLER_29_1004 VPWR VGND sg13g2_decap_8
XFILLER_124_977 VPWR VGND sg13g2_decap_8
X_12145_ _05991_ net1856 fpmul.reg_b_out\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_110_104 VPWR VGND sg13g2_fill_1
XFILLER_111_649 VPWR VGND sg13g2_decap_4
X_12076_ _05922_ _05920_ _05918_ VPWR VGND sg13g2_nand2_1
XFILLER_77_574 VPWR VGND sg13g2_decap_8
X_11027_ VPWR _05006_ _05005_ VGND sg13g2_inv_1
XFILLER_49_265 VPWR VGND sg13g2_decap_4
XFILLER_49_243 VPWR VGND sg13g2_fill_1
XFILLER_38_939 VPWR VGND sg13g2_fill_2
XFILLER_2_56 VPWR VGND sg13g2_decap_8
XFILLER_66_81 VPWR VGND sg13g2_decap_8
XFILLER_64_224 VPWR VGND sg13g2_decap_8
XFILLER_37_438 VPWR VGND sg13g2_decap_8
XFILLER_92_555 VPWR VGND sg13g2_fill_1
XFILLER_92_544 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_29_clk clknet_5_16__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_64_268 VPWR VGND sg13g2_fill_2
XFILLER_52_408 VPWR VGND sg13g2_decap_8
XFILLER_46_950 VPWR VGND sg13g2_decap_8
XFILLER_92_588 VPWR VGND sg13g2_decap_8
XFILLER_75_1013 VPWR VGND sg13g2_fill_1
XFILLER_75_1002 VPWR VGND sg13g2_decap_8
X_12978_ _06746_ _06747_ _06737_ _00894_ VPWR VGND sg13g2_nand3_1
XFILLER_33_600 VPWR VGND sg13g2_decap_8
X_11929_ _05796_ VPWR _00991_ VGND net1879 _05795_ sg13g2_o21ai_1
X_14717_ _00518_ VGND VPWR _01245_ fp16_res_pipe.exp_mant_logic0.a\[4\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
X_14648_ _00449_ VGND VPWR _01176_ fp16_res_pipe.exp_mant_logic0.b\[1\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
XFILLER_60_485 VPWR VGND sg13g2_decap_4
XFILLER_21_839 VPWR VGND sg13g2_decap_8
XFILLER_119_716 VPWR VGND sg13g2_decap_8
XFILLER_9_350 VPWR VGND sg13g2_decap_4
X_14579_ _00380_ VGND VPWR _01111_ fp16_sum_pipe.exp_mant_logic0.b\[6\] clknet_leaf_135_clk
+ sg13g2_dfrbpq_2
XFILLER_9_394 VPWR VGND sg13g2_decap_4
XFILLER_127_771 VPWR VGND sg13g2_decap_8
XFILLER_118_259 VPWR VGND sg13g2_decap_8
XFILLER_115_900 VPWR VGND sg13g2_decap_8
XFILLER_56_0 VPWR VGND sg13g2_decap_8
XFILLER_115_977 VPWR VGND sg13g2_decap_8
XFILLER_87_305 VPWR VGND sg13g2_decap_8
X_07953_ _02227_ fp16_sum_pipe.exp_mant_logic0.b\[8\] VPWR VGND sg13g2_inv_2
X_07884_ _02169_ net1888 acc_sub.x2\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_29_906 VPWR VGND sg13g2_decap_8
X_09623_ net1802 _03740_ VPWR VGND sg13g2_inv_4
XFILLER_28_427 VPWR VGND sg13g2_decap_8
XFILLER_28_449 VPWR VGND sg13g2_fill_1
X_09554_ VGND VPWR _03669_ _02918_ _03671_ _03670_ sg13g2_a21oi_1
XFILLER_70_227 VPWR VGND sg13g2_decap_8
XFILLER_43_419 VPWR VGND sg13g2_decap_4
XFILLER_37_994 VPWR VGND sg13g2_decap_8
XFILLER_36_460 VPWR VGND sg13g2_decap_8
X_08505_ VPWR _02729_ acc_sum.seg_reg1.q\[20\] VGND sg13g2_inv_1
XFILLER_24_622 VPWR VGND sg13g2_fill_1
X_09485_ _03608_ acc_sub.x2\[5\] net1917 VPWR VGND sg13g2_nand2_1
X_08436_ _02670_ _02668_ _02669_ VPWR VGND sg13g2_nand2_1
X_08367_ _02600_ _02609_ _02599_ _02610_ VPWR VGND sg13g2_nand3_1
X_07318_ _01682_ _01541_ _01603_ VPWR VGND sg13g2_nand2b_1
X_08298_ _02545_ net1842 _02408_ fp16_sum_pipe.exp_mant_logic0.b\[6\] _02332_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_125_708 VPWR VGND sg13g2_decap_4
X_07249_ _01487_ _01618_ _01619_ VPWR VGND sg13g2_nand2_1
XFILLER_11_21 VPWR VGND sg13g2_decap_8
XFILLER_127_21 VPWR VGND sg13g2_decap_8
XFILLER_118_782 VPWR VGND sg13g2_decap_8
XFILLER_106_922 VPWR VGND sg13g2_decap_8
XFILLER_3_504 VPWR VGND sg13g2_decap_8
X_10260_ _04330_ VPWR _04331_ VGND _04329_ _04140_ sg13g2_o21ai_1
XFILLER_121_903 VPWR VGND sg13g2_decap_8
XFILLER_11_98 VPWR VGND sg13g2_decap_8
XFILLER_127_98 VPWR VGND sg13g2_decap_8
XFILLER_106_999 VPWR VGND sg13g2_decap_8
XFILLER_105_465 VPWR VGND sg13g2_fill_1
XFILLER_101_660 VPWR VGND sg13g2_decap_8
X_13950_ VPWR _00501_ net97 VGND sg13g2_inv_1
XFILLER_101_671 VPWR VGND sg13g2_fill_2
XFILLER_98_1013 VPWR VGND sg13g2_fill_1
XFILLER_98_1002 VPWR VGND sg13g2_decap_8
XFILLER_86_393 VPWR VGND sg13g2_decap_8
XFILLER_74_533 VPWR VGND sg13g2_fill_2
X_12901_ VPWR _06677_ fpmul.reg_p_out\[6\] VGND sg13g2_inv_1
XFILLER_19_427 VPWR VGND sg13g2_fill_2
XFILLER_100_181 VPWR VGND sg13g2_fill_1
XFILLER_47_758 VPWR VGND sg13g2_decap_8
XFILLER_46_246 VPWR VGND sg13g2_decap_8
X_13881_ VPWR _00432_ net48 VGND sg13g2_inv_1
X_12832_ _06614_ net1716 _00017_ VPWR VGND sg13g2_nand2_1
XFILLER_61_205 VPWR VGND sg13g2_decap_4
XFILLER_46_279 VPWR VGND sg13g2_decap_4
XFILLER_34_419 VPWR VGND sg13g2_fill_2
XFILLER_34_408 VPWR VGND sg13g2_fill_2
XFILLER_15_600 VPWR VGND sg13g2_decap_4
XFILLER_28_994 VPWR VGND sg13g2_decap_8
X_12763_ VGND VPWR net1909 fp16_res_pipe.y\[15\] _06548_ _06547_ sg13g2_a21oi_1
XFILLER_61_238 VPWR VGND sg13g2_decap_8
XFILLER_54_290 VPWR VGND sg13g2_fill_2
XFILLER_36_84 VPWR VGND sg13g2_decap_8
X_14502_ _00303_ VGND VPWR _01038_ fpdiv.reg_b_out\[9\] clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_43_975 VPWR VGND sg13g2_fill_1
XFILLER_15_688 VPWR VGND sg13g2_decap_8
X_11714_ _05618_ _05596_ _05493_ VPWR VGND sg13g2_xnor2_1
X_12694_ VPWR _06503_ _06431_ VGND sg13g2_inv_1
X_14433_ _00234_ VGND VPWR _00972_ fpmul.seg_reg0.q\[18\] clknet_leaf_95_clk sg13g2_dfrbpq_1
XFILLER_11_861 VPWR VGND sg13g2_decap_8
X_11645_ _05550_ _05547_ _05549_ VPWR VGND sg13g2_nand2_1
X_14364_ _00165_ VGND VPWR _00906_ _00017_ clknet_leaf_86_clk sg13g2_dfrbpq_1
XFILLER_7_832 VPWR VGND sg13g2_decap_8
X_11576_ _05480_ VPWR _05481_ VGND net1837 _05424_ sg13g2_o21ai_1
X_13315_ _07023_ _07024_ _07022_ _07025_ VPWR VGND sg13g2_nand3_1
X_14295_ _00096_ VGND VPWR _00839_ acc\[5\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_6_342 VPWR VGND sg13g2_decap_4
X_10527_ net1849 fp16_sum_pipe.add_renorm0.mantisa\[3\] _04568_ VPWR VGND sg13g2_nor2_1
XFILLER_109_793 VPWR VGND sg13g2_decap_8
X_10458_ _04412_ VPWR _04506_ VGND _04500_ _04417_ sg13g2_o21ai_1
XFILLER_124_774 VPWR VGND sg13g2_decap_8
XFILLER_112_936 VPWR VGND sg13g2_decap_8
X_13177_ _06919_ net1715 sipo.word\[11\] VPWR VGND sg13g2_nand2_1
X_10389_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[5\] _04438_ _04439_ VPWR VGND sg13g2_nor2_1
XFILLER_123_273 VPWR VGND sg13g2_decap_8
XFILLER_97_636 VPWR VGND sg13g2_decap_8
X_12128_ _05974_ _05940_ _05973_ VPWR VGND sg13g2_nand2_1
XFILLER_96_157 VPWR VGND sg13g2_decap_8
X_12059_ _05905_ fpmul.reg_b_out\[1\] _05904_ VPWR VGND sg13g2_xnor2_1
XFILLER_77_382 VPWR VGND sg13g2_fill_1
XFILLER_92_341 VPWR VGND sg13g2_fill_2
XFILLER_65_555 VPWR VGND sg13g2_decap_8
XFILLER_37_246 VPWR VGND sg13g2_decap_8
XFILLER_19_950 VPWR VGND sg13g2_decap_8
XFILLER_65_599 VPWR VGND sg13g2_fill_2
XFILLER_53_739 VPWR VGND sg13g2_decap_8
XFILLER_80_536 VPWR VGND sg13g2_decap_8
XFILLER_45_290 VPWR VGND sg13g2_fill_1
XFILLER_34_975 VPWR VGND sg13g2_decap_8
X_09270_ fp16_res_pipe.op_sign_logic0.mantisa_b\[4\] _03423_ _03424_ VPWR VGND sg13g2_nor2_1
XFILLER_20_113 VPWR VGND sg13g2_decap_8
XFILLER_21_636 VPWR VGND sg13g2_decap_8
XFILLER_33_485 VPWR VGND sg13g2_fill_2
X_08152_ _02406_ _02411_ _02412_ VPWR VGND sg13g2_nor2_1
XFILLER_20_179 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_9_clk clknet_5_4__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_08083_ _02349_ _02347_ VPWR VGND sg13g2_inv_2
Xclkbuf_5_15__f_clk clknet_4_7_0_clk clknet_5_15__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_127_590 VPWR VGND sg13g2_decap_8
XFILLER_115_774 VPWR VGND sg13g2_decap_8
XFILLER_103_925 VPWR VGND sg13g2_decap_8
X_08985_ VPWR _03171_ _03170_ VGND sg13g2_inv_1
XFILLER_114_284 VPWR VGND sg13g2_decap_8
XFILLER_87_146 VPWR VGND sg13g2_decap_8
XFILLER_69_850 VPWR VGND sg13g2_decap_4
X_07936_ fp16_sum_pipe.exp_mant_logic0.a\[9\] _02210_ _02211_ VPWR VGND sg13g2_nor2_1
XFILLER_84_831 VPWR VGND sg13g2_fill_2
XFILLER_68_360 VPWR VGND sg13g2_decap_8
XFILLER_56_511 VPWR VGND sg13g2_decap_4
XFILLER_29_725 VPWR VGND sg13g2_fill_2
X_07867_ _02160_ VPWR _01410_ VGND acc_sub.reg1en.q\[0\] _01545_ sg13g2_o21ai_1
XFILLER_84_853 VPWR VGND sg13g2_decap_8
XFILLER_56_555 VPWR VGND sg13g2_decap_4
XFILLER_56_544 VPWR VGND sg13g2_decap_8
XFILLER_44_706 VPWR VGND sg13g2_fill_1
XFILLER_28_246 VPWR VGND sg13g2_fill_2
XFILLER_113_56 VPWR VGND sg13g2_decap_8
X_09606_ net1805 acc_sum.add_renorm0.mantisa\[10\] _03723_ VPWR VGND sg13g2_nor2_2
X_07798_ _02096_ _02024_ _02097_ VPWR VGND sg13g2_nor2_1
XFILLER_71_514 VPWR VGND sg13g2_decap_8
XFILLER_56_588 VPWR VGND sg13g2_decap_8
X_09537_ VPWR _03654_ _03652_ VGND sg13g2_inv_1
XFILLER_25_931 VPWR VGND sg13g2_decap_8
XFILLER_40_901 VPWR VGND sg13g2_fill_2
XFILLER_106_1006 VPWR VGND sg13g2_decap_8
XFILLER_51_271 VPWR VGND sg13g2_fill_2
X_09468_ _03596_ VPWR _01252_ VGND net1914 _03595_ sg13g2_o21ai_1
X_08419_ net1707 fpdiv.divider0.en_r VPWR VGND sg13g2_inv_4
XFILLER_40_978 VPWR VGND sg13g2_decap_8
XFILLER_8_607 VPWR VGND sg13g2_decap_8
X_09399_ _03544_ VPWR _03545_ VGND _03425_ _03543_ sg13g2_o21ai_1
X_11430_ VPWR _05363_ fpdiv.reg_a_out\[11\] VGND sg13g2_inv_1
XFILLER_22_42 VPWR VGND sg13g2_decap_8
X_11361_ _05310_ _05312_ _05313_ VPWR VGND sg13g2_nor2_1
X_13100_ _06859_ VPWR _00884_ VGND net1862 _06677_ sg13g2_o21ai_1
X_10312_ _04373_ VPWR _01185_ VGND net1914 _04018_ sg13g2_o21ai_1
XFILLER_3_301 VPWR VGND sg13g2_decap_4
X_14080_ VPWR _00631_ net138 VGND sg13g2_inv_1
X_11292_ _05248_ _05249_ _05250_ _05252_ VGND VPWR _05251_ sg13g2_nor4_2
XFILLER_4_846 VPWR VGND sg13g2_decap_8
XFILLER_106_774 VPWR VGND sg13g2_fill_2
XFILLER_79_603 VPWR VGND sg13g2_fill_1
X_13031_ _06799_ _06796_ _06797_ _06798_ VPWR VGND sg13g2_and3_1
XFILLER_3_378 VPWR VGND sg13g2_decap_8
X_10243_ _04313_ _04314_ _04315_ VPWR VGND sg13g2_and2_1
XFILLER_120_210 VPWR VGND sg13g2_decap_8
XFILLER_79_647 VPWR VGND sg13g2_fill_2
X_10174_ _04254_ net1764 fp16_res_pipe.op_sign_logic0.mantisa_a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_121_777 VPWR VGND sg13g2_decap_8
XFILLER_78_168 VPWR VGND sg13g2_decap_4
XFILLER_120_287 VPWR VGND sg13g2_fill_1
XFILLER_94_628 VPWR VGND sg13g2_decap_8
XFILLER_59_382 VPWR VGND sg13g2_fill_1
XFILLER_59_371 VPWR VGND sg13g2_fill_1
XFILLER_19_213 VPWR VGND sg13g2_fill_2
XFILLER_75_842 VPWR VGND sg13g2_decap_4
XFILLER_47_61 VPWR VGND sg13g2_decap_8
X_13933_ VPWR _00484_ net6 VGND sg13g2_inv_1
XFILLER_74_374 VPWR VGND sg13g2_fill_1
XFILLER_74_363 VPWR VGND sg13g2_decap_8
XFILLER_47_566 VPWR VGND sg13g2_decap_8
X_13864_ VPWR _00415_ net52 VGND sg13g2_inv_1
XFILLER_35_728 VPWR VGND sg13g2_decap_8
XFILLER_34_216 VPWR VGND sg13g2_fill_1
X_12815_ _06598_ _06594_ _06597_ _06593_ net1941 VPWR VGND sg13g2_a22oi_1
XFILLER_16_931 VPWR VGND sg13g2_decap_8
XFILLER_90_889 VPWR VGND sg13g2_decap_8
XFILLER_90_878 VPWR VGND sg13g2_fill_1
X_13795_ VPWR _00346_ net20 VGND sg13g2_inv_1
XFILLER_43_750 VPWR VGND sg13g2_decap_8
XFILLER_27_290 VPWR VGND sg13g2_decap_8
XFILLER_97_7 VPWR VGND sg13g2_fill_2
X_12746_ fpmul.reg_b_out\[11\] fp16_res_pipe.x2\[11\] net1952 _00921_ VPWR VGND sg13g2_mux2_1
XFILLER_30_411 VPWR VGND sg13g2_decap_8
X_12677_ VPWR _06490_ _06360_ VGND sg13g2_inv_1
XFILLER_31_956 VPWR VGND sg13g2_decap_8
X_14416_ _00217_ VGND VPWR _00955_ fpmul.reg_a_out\[13\] clknet_leaf_125_clk sg13g2_dfrbpq_2
X_11628_ _05533_ _05532_ _05520_ VPWR VGND sg13g2_nand2_1
X_14347_ _00148_ VGND VPWR _00889_ fpmul.reg_p_out\[11\] clknet_leaf_89_clk sg13g2_dfrbpq_1
XFILLER_8_77 VPWR VGND sg13g2_decap_8
XFILLER_6_161 VPWR VGND sg13g2_decap_8
X_11559_ VPWR _05464_ _05455_ VGND sg13g2_inv_1
XFILLER_116_549 VPWR VGND sg13g2_decap_8
X_14278_ _00079_ VGND VPWR _00829_ fp16_res_pipe.x2\[11\] clknet_leaf_130_clk sg13g2_dfrbpq_2
XFILLER_98_912 VPWR VGND sg13g2_fill_2
X_13229_ acc_sum.reg4en.q\[0\] _02573_ _06954_ VPWR VGND sg13g2_nor2_1
XFILLER_98_967 VPWR VGND sg13g2_decap_8
XFILLER_97_411 VPWR VGND sg13g2_decap_8
XFILLER_111_254 VPWR VGND sg13g2_decap_8
XFILLER_97_499 VPWR VGND sg13g2_decap_8
X_08770_ _02960_ acc\[2\] net1896 VPWR VGND sg13g2_nand2_1
X_07721_ _02028_ _02021_ _02027_ VPWR VGND sg13g2_nand2_1
XFILLER_84_138 VPWR VGND sg13g2_fill_1
XFILLER_77_190 VPWR VGND sg13g2_fill_1
XFILLER_38_544 VPWR VGND sg13g2_decap_8
XFILLER_19_0 VPWR VGND sg13g2_decap_8
X_07652_ _01964_ net1641 _01963_ VPWR VGND sg13g2_nand2_1
XFILLER_38_599 VPWR VGND sg13g2_fill_2
X_07583_ VGND VPWR _01893_ _01792_ _01897_ _01896_ sg13g2_a21oi_1
XFILLER_53_547 VPWR VGND sg13g2_decap_8
XFILLER_25_216 VPWR VGND sg13g2_decap_8
XFILLER_25_227 VPWR VGND sg13g2_fill_2
X_09322_ _03475_ _03474_ _03437_ VPWR VGND sg13g2_nand2_1
XFILLER_22_912 VPWR VGND sg13g2_decap_8
XFILLER_61_580 VPWR VGND sg13g2_decap_4
XFILLER_40_219 VPWR VGND sg13g2_decap_8
XFILLER_21_411 VPWR VGND sg13g2_decap_4
X_09253_ _03404_ _03406_ _03407_ VPWR VGND sg13g2_nor2_2
XFILLER_21_433 VPWR VGND sg13g2_decap_8
XFILLER_119_321 VPWR VGND sg13g2_decap_8
X_09184_ _03346_ acc_sub.x2\[6\] net1905 VPWR VGND sg13g2_nand2_1
X_08204_ _02460_ fp16_sum_pipe.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_inv_2
XFILLER_21_477 VPWR VGND sg13g2_decap_8
XFILLER_22_989 VPWR VGND sg13g2_decap_8
X_08135_ _02307_ _02328_ _02396_ VPWR VGND _02336_ sg13g2_nand3b_1
XFILLER_119_398 VPWR VGND sg13g2_fill_2
X_08066_ _02305_ _02331_ _02332_ VPWR VGND sg13g2_nor2b_2
XFILLER_115_560 VPWR VGND sg13g2_decap_4
XFILLER_108_67 VPWR VGND sg13g2_decap_8
Xplace1851 fpdiv.div_out\[11\] net1851 VPWR VGND sg13g2_buf_2
XFILLER_68_16 VPWR VGND sg13g2_decap_4
Xplace1862 fpmul.reg2en.q\[0\] net1862 VPWR VGND sg13g2_buf_2
Xplace1840 fp16_sum_pipe.add_renorm0.mantisa\[11\] net1840 VPWR VGND sg13g2_buf_2
XFILLER_115_593 VPWR VGND sg13g2_decap_8
Xplace1895 net1893 net1895 VPWR VGND sg13g2_buf_2
XFILLER_88_411 VPWR VGND sg13g2_decap_8
Xplace1873 fpmul.reg1en.q\[0\] net1873 VPWR VGND sg13g2_buf_2
Xplace1884 net1883 net1884 VPWR VGND sg13g2_buf_2
XFILLER_0_337 VPWR VGND sg13g2_decap_8
X_08968_ _03154_ acc_sub.add_renorm0.exp\[3\] _03139_ VPWR VGND sg13g2_xnor2_1
XFILLER_102_276 VPWR VGND sg13g2_fill_2
XFILLER_88_499 VPWR VGND sg13g2_decap_8
XFILLER_76_639 VPWR VGND sg13g2_decap_8
XFILLER_75_127 VPWR VGND sg13g2_decap_4
X_08899_ _03085_ VPWR _03086_ VGND _03082_ _03084_ sg13g2_o21ai_1
XFILLER_124_77 VPWR VGND sg13g2_decap_8
XFILLER_29_555 VPWR VGND sg13g2_decap_8
X_07919_ _02194_ fp16_sum_pipe.exp_mant_logic0.b\[11\] VPWR VGND sg13g2_inv_2
XFILLER_84_672 VPWR VGND sg13g2_decap_8
XFILLER_17_717 VPWR VGND sg13g2_decap_8
X_10930_ net1771 VPWR _04938_ VGND _04937_ _04924_ sg13g2_o21ai_1
XFILLER_72_834 VPWR VGND sg13g2_decap_8
XFILLER_17_42 VPWR VGND sg13g2_decap_8
XFILLER_17_739 VPWR VGND sg13g2_decap_4
XFILLER_29_599 VPWR VGND sg13g2_decap_4
XFILLER_72_889 VPWR VGND sg13g2_decap_8
XFILLER_72_867 VPWR VGND sg13g2_decap_4
X_12600_ _06395_ _06407_ _06416_ VPWR VGND sg13g2_xor2_1
X_10861_ VGND VPWR _04800_ net1824 _04873_ _04872_ sg13g2_a21oi_1
X_13580_ VPWR _00131_ net120 VGND sg13g2_inv_1
XFILLER_40_720 VPWR VGND sg13g2_decap_8
XFILLER_13_912 VPWR VGND sg13g2_decap_8
X_10792_ _03584_ VPWR _04804_ VGND _03586_ _04803_ sg13g2_o21ai_1
X_12531_ _06351_ VPWR _00944_ VGND net1954 _05913_ sg13g2_o21ai_1
XFILLER_8_404 VPWR VGND sg13g2_decap_8
XFILLER_9_927 VPWR VGND sg13g2_decap_8
X_12462_ VPWR _06304_ fpmul.seg_reg0.q\[11\] VGND sg13g2_inv_1
XFILLER_13_989 VPWR VGND sg13g2_decap_8
XFILLER_33_63 VPWR VGND sg13g2_decap_8
XFILLER_123_0 VPWR VGND sg13g2_decap_8
X_14201_ VPWR _00752_ net105 VGND sg13g2_inv_1
X_11413_ _05352_ VPWR _01063_ VGND _05350_ fpdiv.divider0.en_r sg13g2_o21ai_1
X_12393_ _06239_ _06220_ _06221_ VPWR VGND sg13g2_xnor2_1
XFILLER_126_869 VPWR VGND sg13g2_decap_8
X_14132_ VPWR _00683_ net102 VGND sg13g2_inv_1
X_11344_ _05297_ net1654 acc_sum.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
X_14063_ VPWR _00614_ net94 VGND sg13g2_inv_1
X_11275_ _05237_ net1808 _05227_ net1809 _05211_ VPWR VGND sg13g2_a22oi_1
X_13014_ net1853 fpmul.seg_reg0.q\[9\] _06782_ VPWR VGND sg13g2_nor2_1
XFILLER_3_175 VPWR VGND sg13g2_decap_8
X_10226_ _04298_ net1703 _04299_ VPWR VGND sg13g2_nor2_1
XFILLER_121_530 VPWR VGND sg13g2_decap_8
XFILLER_94_414 VPWR VGND sg13g2_decap_4
XFILLER_94_403 VPWR VGND sg13g2_fill_1
XFILLER_79_488 VPWR VGND sg13g2_decap_8
X_10157_ _04237_ VPWR _04238_ VGND _03617_ _04124_ sg13g2_o21ai_1
X_14965_ _00766_ VGND VPWR _01485_ acc_sub.add_renorm0.mantisa\[9\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_2
XFILLER_12_7 VPWR VGND sg13g2_decap_8
X_10088_ _04173_ _04076_ fp16_res_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_81_108 VPWR VGND sg13g2_decap_4
X_13916_ VPWR _00467_ net8 VGND sg13g2_inv_1
X_14896_ _00697_ VGND VPWR _01416_ acc_sub.op_sign_logic0.mantisa_b\[6\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_1
XFILLER_90_631 VPWR VGND sg13g2_decap_8
XFILLER_62_322 VPWR VGND sg13g2_fill_2
XFILLER_35_525 VPWR VGND sg13g2_decap_8
XFILLER_74_81 VPWR VGND sg13g2_decap_4
XFILLER_63_889 VPWR VGND sg13g2_decap_8
X_13847_ VPWR _00398_ net29 VGND sg13g2_inv_1
X_13778_ VPWR _00329_ net125 VGND sg13g2_inv_1
XFILLER_16_783 VPWR VGND sg13g2_decap_8
X_12729_ VPWR _06533_ div_result\[2\] VGND sg13g2_inv_1
XFILLER_30_285 VPWR VGND sg13g2_fill_1
XFILLER_30_296 VPWR VGND sg13g2_fill_2
XFILLER_8_993 VPWR VGND sg13g2_decap_8
XFILLER_117_858 VPWR VGND sg13g2_decap_8
XFILLER_116_335 VPWR VGND sg13g2_fill_1
XFILLER_7_470 VPWR VGND sg13g2_decap_8
X_09940_ _04035_ VPWR _04036_ VGND _04013_ _04010_ sg13g2_o21ai_1
XFILLER_124_390 VPWR VGND sg13g2_fill_1
X_09871_ _03977_ _03631_ _03666_ _03635_ _03630_ VPWR VGND sg13g2_a22oi_1
XFILLER_98_775 VPWR VGND sg13g2_decap_8
XFILLER_97_241 VPWR VGND sg13g2_fill_1
X_08822_ net1704 _03009_ VPWR VGND sg13g2_inv_4
XFILLER_112_596 VPWR VGND sg13g2_fill_2
XFILLER_86_959 VPWR VGND sg13g2_decap_8
XFILLER_85_458 VPWR VGND sg13g2_fill_1
XFILLER_85_436 VPWR VGND sg13g2_fill_2
X_08753_ _02948_ VPWR _01319_ VGND net1900 _02947_ sg13g2_o21ai_1
X_07704_ _02012_ _02011_ _01944_ VPWR VGND sg13g2_nand2_1
XFILLER_39_875 VPWR VGND sg13g2_decap_8
XFILLER_38_352 VPWR VGND sg13g2_fill_1
X_08684_ net1817 acc_sum.add_renorm0.mantisa\[4\] _02900_ VPWR VGND sg13g2_nor2_1
XFILLER_93_491 VPWR VGND sg13g2_fill_1
X_07635_ _01430_ _01946_ _01948_ VPWR VGND sg13g2_nand2_1
XFILLER_81_664 VPWR VGND sg13g2_fill_1
XFILLER_65_193 VPWR VGND sg13g2_decap_8
XFILLER_110_35 VPWR VGND sg13g2_decap_8
X_07566_ VPWR _01880_ _01812_ VGND sg13g2_inv_1
XFILLER_80_185 VPWR VGND sg13g2_decap_4
XFILLER_41_528 VPWR VGND sg13g2_fill_1
XFILLER_13_208 VPWR VGND sg13g2_decap_4
X_09305_ _03458_ VPWR _01277_ VGND net1833 _03367_ sg13g2_o21ai_1
X_07497_ _01811_ _01819_ _01820_ VPWR VGND sg13g2_nor2_1
X_09236_ _03383_ _03389_ _03390_ VPWR VGND sg13g2_nor2_1
XFILLER_10_926 VPWR VGND sg13g2_decap_8
XFILLER_103_1009 VPWR VGND sg13g2_decap_4
XFILLER_119_140 VPWR VGND sg13g2_decap_8
X_09167_ _03334_ VPWR _01291_ VGND net1904 _03333_ sg13g2_o21ai_1
XFILLER_5_429 VPWR VGND sg13g2_decap_8
XFILLER_5_407 VPWR VGND sg13g2_decap_4
XFILLER_119_77 VPWR VGND sg13g2_decap_8
X_09098_ VGND VPWR net1786 _03280_ _03281_ _03136_ sg13g2_a21oi_1
X_08118_ _02380_ net1657 VPWR VGND sg13g2_inv_2
XFILLER_123_806 VPWR VGND sg13g2_decap_8
X_08049_ _02315_ _02311_ _02314_ VPWR VGND sg13g2_nand2_1
XFILLER_116_891 VPWR VGND sg13g2_decap_8
X_11060_ VPWR _05038_ _04999_ VGND sg13g2_inv_1
Xplace1681 _05049_ net1681 VPWR VGND sg13g2_buf_2
XFILLER_0_112 VPWR VGND sg13g2_decap_8
Xplace1670 _04530_ net1670 VPWR VGND sg13g2_buf_2
XFILLER_115_390 VPWR VGND sg13g2_decap_4
XFILLER_88_230 VPWR VGND sg13g2_decap_8
X_10011_ _04098_ VPWR _04099_ VGND _04077_ _04050_ sg13g2_o21ai_1
Xplace1692 _02244_ net1692 VPWR VGND sg13g2_buf_2
XFILLER_103_574 VPWR VGND sg13g2_fill_1
XFILLER_77_948 VPWR VGND sg13g2_decap_8
XFILLER_77_937 VPWR VGND sg13g2_fill_1
XFILLER_76_403 VPWR VGND sg13g2_fill_1
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_103_596 VPWR VGND sg13g2_decap_4
XFILLER_76_458 VPWR VGND sg13g2_decap_4
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_91_428 VPWR VGND sg13g2_decap_4
XFILLER_91_406 VPWR VGND sg13g2_fill_1
XFILLER_57_661 VPWR VGND sg13g2_fill_1
XFILLER_45_812 VPWR VGND sg13g2_decap_8
X_14750_ _00551_ VGND VPWR _01278_ fp16_res_pipe.seg_reg1.q\[21\] clknet_leaf_139_clk
+ sg13g2_dfrbpq_2
XFILLER_28_63 VPWR VGND sg13g2_decap_8
XFILLER_85_992 VPWR VGND sg13g2_decap_8
XFILLER_84_480 VPWR VGND sg13g2_decap_8
XFILLER_56_182 VPWR VGND sg13g2_decap_8
X_11962_ _05818_ VPWR _00980_ VGND net1884 _05817_ sg13g2_o21ai_1
XFILLER_45_823 VPWR VGND sg13g2_fill_1
X_13701_ VPWR _00252_ net54 VGND sg13g2_inv_1
XFILLER_44_300 VPWR VGND sg13g2_decap_8
XFILLER_29_385 VPWR VGND sg13g2_fill_1
X_11893_ fpmul.result\[15\] net1876 _05778_ VPWR VGND sg13g2_nor2_1
X_14681_ _00482_ VGND VPWR _01209_ fp16_res_pipe.op_sign_logic0.mantisa_a\[7\] clknet_leaf_143_clk
+ sg13g2_dfrbpq_2
X_10913_ _04743_ VPWR _04922_ VGND _04829_ _04921_ sg13g2_o21ai_1
XFILLER_71_185 VPWR VGND sg13g2_decap_8
X_13632_ VPWR _00183_ net50 VGND sg13g2_inv_1
X_10844_ _04856_ _04834_ _04855_ VPWR VGND sg13g2_nand2_1
X_13563_ VPWR _00114_ net82 VGND sg13g2_inv_1
XFILLER_44_84 VPWR VGND sg13g2_decap_8
X_12514_ VGND VPWR _06341_ net1953 _00952_ _06342_ sg13g2_a21oi_1
XFILLER_9_724 VPWR VGND sg13g2_fill_2
XFILLER_12_252 VPWR VGND sg13g2_decap_8
XFILLER_13_786 VPWR VGND sg13g2_decap_4
X_13494_ VPWR _00045_ net35 VGND sg13g2_inv_1
XFILLER_8_234 VPWR VGND sg13g2_fill_1
XFILLER_9_757 VPWR VGND sg13g2_decap_8
XFILLER_126_611 VPWR VGND sg13g2_decap_8
X_12445_ _06285_ _06290_ _06289_ _06291_ VPWR VGND sg13g2_nand3_1
XFILLER_8_256 VPWR VGND sg13g2_decap_4
XFILLER_126_633 VPWR VGND sg13g2_fill_1
X_12376_ _06220_ _06221_ _06222_ VPWR VGND sg13g2_nor2_1
XFILLER_5_941 VPWR VGND sg13g2_decap_8
XFILLER_125_154 VPWR VGND sg13g2_decap_8
X_11327_ _03349_ _05173_ _05282_ VPWR VGND sg13g2_nor2_1
X_14115_ VPWR _00666_ net52 VGND sg13g2_inv_1
XFILLER_114_839 VPWR VGND sg13g2_decap_8
XFILLER_113_327 VPWR VGND sg13g2_fill_1
XFILLER_5_56 VPWR VGND sg13g2_decap_8
XFILLER_4_462 VPWR VGND sg13g2_decap_8
XFILLER_122_861 VPWR VGND sg13g2_decap_8
XFILLER_79_230 VPWR VGND sg13g2_decap_8
X_14046_ VPWR _00597_ net86 VGND sg13g2_inv_1
X_11258_ _05220_ VPWR _05221_ VGND _02959_ _05143_ sg13g2_o21ai_1
XFILLER_95_734 VPWR VGND sg13g2_fill_1
X_11189_ _05158_ net1635 _05157_ VPWR VGND sg13g2_nand2_1
XFILLER_39_105 VPWR VGND sg13g2_decap_8
X_10209_ _04284_ net1644 net1830 VPWR VGND sg13g2_nand2_1
XFILLER_121_393 VPWR VGND sg13g2_fill_2
XFILLER_95_745 VPWR VGND sg13g2_decap_8
XFILLER_94_233 VPWR VGND sg13g2_decap_8
XFILLER_95_778 VPWR VGND sg13g2_fill_2
XFILLER_83_918 VPWR VGND sg13g2_decap_8
XFILLER_76_981 VPWR VGND sg13g2_fill_2
X_14948_ _00749_ VGND VPWR _01468_ acc_sub.add_renorm0.exp\[0\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_2
XFILLER_91_940 VPWR VGND sg13g2_decap_8
XFILLER_82_439 VPWR VGND sg13g2_decap_4
XFILLER_78_1011 VPWR VGND sg13g2_fill_2
XFILLER_63_620 VPWR VGND sg13g2_fill_1
XFILLER_48_694 VPWR VGND sg13g2_decap_4
XFILLER_47_171 VPWR VGND sg13g2_fill_2
X_14879_ _00680_ VGND VPWR _01399_ acc_sub.exp_mant_logic0.b\[5\] clknet_leaf_58_clk
+ sg13g2_dfrbpq_1
XFILLER_126_1009 VPWR VGND sg13g2_decap_4
X_07420_ VPWR _01755_ fpdiv.reg1en.q\[0\] VGND sg13g2_inv_1
XFILLER_35_366 VPWR VGND sg13g2_decap_8
X_07351_ _01710_ net1799 acc_sub.seg_reg0.q\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_16_580 VPWR VGND sg13g2_decap_8
XFILLER_86_0 VPWR VGND sg13g2_decap_8
XFILLER_31_550 VPWR VGND sg13g2_fill_2
X_07282_ net1783 _01648_ _01649_ _01650_ VPWR VGND sg13g2_nor3_1
XFILLER_31_583 VPWR VGND sg13g2_fill_1
X_09021_ _03207_ _03205_ _03206_ VPWR VGND sg13g2_nand2_1
XFILLER_116_110 VPWR VGND sg13g2_decap_8
XFILLER_117_655 VPWR VGND sg13g2_decap_8
XFILLER_116_187 VPWR VGND sg13g2_decap_8
XFILLER_105_839 VPWR VGND sg13g2_fill_2
X_09923_ _04020_ _03597_ fp16_res_pipe.exp_mant_logic0.b\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_113_872 VPWR VGND sg13g2_decap_8
X_09854_ _03964_ _03961_ _03963_ _03958_ net1769 VPWR VGND sg13g2_a22oi_1
X_08805_ _02992_ _02976_ acc_sub.add_renorm0.mantisa\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_112_382 VPWR VGND sg13g2_fill_2
XFILLER_100_533 VPWR VGND sg13g2_decap_8
XFILLER_86_745 VPWR VGND sg13g2_fill_1
XFILLER_105_79 VPWR VGND sg13g2_fill_2
X_09785_ _03783_ _03899_ _03896_ _03900_ VPWR VGND sg13g2_nand3_1
XFILLER_65_28 VPWR VGND sg13g2_decap_8
XFILLER_22_1010 VPWR VGND sg13g2_decap_4
XFILLER_100_588 VPWR VGND sg13g2_decap_8
XFILLER_82_940 VPWR VGND sg13g2_decap_8
XFILLER_73_439 VPWR VGND sg13g2_decap_8
XFILLER_67_992 VPWR VGND sg13g2_fill_2
X_08736_ _02937_ acc_sum.exp_mant_logic0.a\[13\] VPWR VGND sg13g2_inv_2
XFILLER_45_119 VPWR VGND sg13g2_decap_8
XFILLER_26_300 VPWR VGND sg13g2_fill_2
X_08667_ _02885_ net1668 _02785_ VPWR VGND sg13g2_nand2b_1
XFILLER_121_56 VPWR VGND sg13g2_decap_8
X_07618_ _01871_ _01923_ _01931_ _01932_ VPWR VGND sg13g2_nor3_1
XFILLER_81_16 VPWR VGND sg13g2_decap_8
XFILLER_53_163 VPWR VGND sg13g2_decap_8
X_08598_ VGND VPWR _02816_ _02818_ _02821_ _02820_ sg13g2_a21oi_1
XFILLER_81_494 VPWR VGND sg13g2_fill_1
X_07549_ _01745_ _01751_ _01743_ _01864_ VPWR VGND sg13g2_nand3_1
XFILLER_14_21 VPWR VGND sg13g2_decap_8
X_10560_ _04592_ fp16_sum_pipe.seg_reg0.q\[24\] net1845 VPWR VGND sg13g2_nand2_1
XFILLER_127_419 VPWR VGND sg13g2_decap_8
X_10491_ VGND VPWR _04447_ _04408_ _04536_ _04407_ sg13g2_a21oi_1
X_09219_ fp16_res_pipe.op_sign_logic0.mantisa_b\[9\] _03372_ _03373_ VPWR VGND sg13g2_nor2_1
X_12230_ _06075_ _06071_ _06076_ VPWR VGND sg13g2_xor2_1
XFILLER_30_42 VPWR VGND sg13g2_decap_8
XFILLER_123_614 VPWR VGND sg13g2_decap_4
X_12161_ _06007_ _06006_ _05985_ VPWR VGND sg13g2_nand2_1
XFILLER_2_933 VPWR VGND sg13g2_decap_8
XFILLER_107_198 VPWR VGND sg13g2_decap_8
X_11112_ _05080_ _05081_ _05082_ VPWR VGND sg13g2_nor2b_1
X_12092_ _05938_ _05933_ _05937_ VPWR VGND sg13g2_nand2_1
XFILLER_1_443 VPWR VGND sg13g2_decap_8
XFILLER_122_168 VPWR VGND sg13g2_decap_8
X_11043_ acc_sum.exp_mant_logic0.b\[7\] _02949_ _05022_ VPWR VGND sg13g2_nor2_2
XFILLER_77_701 VPWR VGND sg13g2_decap_4
XFILLER_49_403 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_92_726 VPWR VGND sg13g2_decap_8
XFILLER_92_715 VPWR VGND sg13g2_decap_8
X_14802_ _00603_ VGND VPWR _01326_ acc_sum.exp_mant_logic0.a\[15\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
Xclkbuf_4_3_0_clk clknet_0_clk clknet_4_3_0_clk VPWR VGND sg13g2_buf_8
XFILLER_91_225 VPWR VGND sg13g2_decap_8
XFILLER_76_299 VPWR VGND sg13g2_fill_1
XFILLER_76_288 VPWR VGND sg13g2_decap_8
X_12994_ _06751_ fpmul.seg_reg0.q\[18\] _06762_ VPWR VGND sg13g2_xor2_1
XFILLER_36_119 VPWR VGND sg13g2_fill_2
XFILLER_73_973 VPWR VGND sg13g2_decap_8
X_11945_ VPWR _05807_ fpmul.seg_reg0.q\[31\] VGND sg13g2_inv_1
XFILLER_45_664 VPWR VGND sg13g2_decap_8
XFILLER_18_878 VPWR VGND sg13g2_decap_8
X_14733_ _00534_ VGND VPWR _01261_ fp16_res_pipe.add_renorm0.exp\[4\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_1
XFILLER_60_601 VPWR VGND sg13g2_fill_2
XFILLER_55_94 VPWR VGND sg13g2_decap_8
X_14664_ _00465_ VGND VPWR _01192_ fp16_res_pipe.op_sign_logic0.mantisa_b\[1\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_1
X_13615_ VPWR _00166_ net112 VGND sg13g2_inv_1
X_11876_ _05765_ VPWR _01013_ VGND net1850 _05764_ sg13g2_o21ai_1
XFILLER_60_678 VPWR VGND sg13g2_fill_1
X_14595_ _00396_ VGND VPWR _01127_ fp16_res_pipe.y\[6\] clknet_leaf_128_clk sg13g2_dfrbpq_1
XFILLER_41_870 VPWR VGND sg13g2_fill_2
XFILLER_13_561 VPWR VGND sg13g2_decap_8
X_10827_ _04839_ _04838_ _04667_ VPWR VGND sg13g2_nand2_1
X_13546_ VPWR _00097_ net101 VGND sg13g2_inv_1
X_10758_ _04771_ _04770_ fp16_res_pipe.reg3en.q\[0\] VPWR VGND sg13g2_nand2_2
XFILLER_71_93 VPWR VGND sg13g2_decap_8
X_13477_ VPWR _00028_ net26 VGND sg13g2_inv_1
XFILLER_9_576 VPWR VGND sg13g2_fill_2
XFILLER_127_953 VPWR VGND sg13g2_decap_8
X_12428_ _06258_ _06259_ _06274_ VPWR VGND sg13g2_nor2_1
X_10689_ _04701_ VPWR _04702_ VGND net1822 _04691_ sg13g2_o21ai_1
XFILLER_126_496 VPWR VGND sg13g2_fill_1
XFILLER_114_636 VPWR VGND sg13g2_decap_8
XFILLER_99_303 VPWR VGND sg13g2_decap_4
X_12359_ _06172_ _06198_ _06200_ _06205_ VPWR VGND sg13g2_nand3_1
XFILLER_113_135 VPWR VGND sg13g2_fill_1
X_14029_ VPWR _00580_ net99 VGND sg13g2_inv_1
XFILLER_68_723 VPWR VGND sg13g2_decap_8
XFILLER_68_756 VPWR VGND sg13g2_decap_8
XFILLER_110_864 VPWR VGND sg13g2_decap_8
XFILLER_67_266 VPWR VGND sg13g2_decap_8
XFILLER_67_244 VPWR VGND sg13g2_fill_2
X_09570_ VPWR _03687_ _03680_ VGND sg13g2_inv_1
XFILLER_95_586 VPWR VGND sg13g2_decap_8
XFILLER_49_981 VPWR VGND sg13g2_decap_8
XFILLER_48_480 VPWR VGND sg13g2_fill_1
XFILLER_27_119 VPWR VGND sg13g2_decap_4
X_08521_ _02738_ _02744_ _02745_ VPWR VGND sg13g2_nor2_1
XFILLER_82_258 VPWR VGND sg13g2_fill_1
X_08452_ _02685_ VPWR _02686_ VGND fpdiv.divider0.remainder_reg\[11\] _02683_ sg13g2_o21ai_1
XFILLER_91_792 VPWR VGND sg13g2_fill_1
XFILLER_63_472 VPWR VGND sg13g2_fill_2
XFILLER_36_697 VPWR VGND sg13g2_decap_8
X_07403_ _01744_ net1887 acc\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_50_133 VPWR VGND sg13g2_decap_8
X_08383_ _02622_ _07114_ fp16_sum_pipe.reg4en.q\[0\] VPWR VGND sg13g2_nand2b_1
XFILLER_11_509 VPWR VGND sg13g2_decap_8
X_07334_ _01636_ VPWR _01696_ VGND _01564_ _01694_ sg13g2_o21ai_1
XFILLER_31_380 VPWR VGND sg13g2_decap_8
X_07265_ VPWR _01635_ _01495_ VGND sg13g2_inv_1
X_09004_ _03153_ _03189_ _03190_ VPWR VGND sg13g2_nor2_1
X_07196_ VPWR _01568_ _01555_ VGND sg13g2_inv_1
XFILLER_118_964 VPWR VGND sg13g2_decap_8
XFILLER_117_474 VPWR VGND sg13g2_decap_8
XFILLER_116_12 VPWR VGND sg13g2_decap_8
X_09906_ VPWR _04003_ _04002_ VGND sg13g2_inv_1
XFILLER_116_89 VPWR VGND sg13g2_decap_8
XFILLER_101_842 VPWR VGND sg13g2_decap_8
XFILLER_59_734 VPWR VGND sg13g2_fill_2
X_09837_ _03628_ _03851_ _03948_ VPWR VGND sg13g2_nor2_1
XFILLER_47_918 VPWR VGND sg13g2_fill_1
X_09768_ _03663_ VPWR _03884_ VGND _03865_ _03883_ sg13g2_o21ai_1
XFILLER_100_396 VPWR VGND sg13g2_fill_1
XFILLER_100_385 VPWR VGND sg13g2_decap_8
XFILLER_18_108 VPWR VGND sg13g2_decap_8
XFILLER_18_119 VPWR VGND sg13g2_fill_2
X_08719_ VPWR _02926_ acc_sum.add_renorm0.exp\[3\] VGND sg13g2_inv_1
XFILLER_73_236 VPWR VGND sg13g2_fill_1
X_09699_ _03815_ acc_sum.add_renorm0.exp\[4\] _03789_ VPWR VGND sg13g2_xnor2_1
XFILLER_70_921 VPWR VGND sg13g2_decap_4
X_11730_ _05634_ _05633_ _05592_ VPWR VGND sg13g2_nand2_1
XFILLER_25_42 VPWR VGND sg13g2_decap_8
XFILLER_42_667 VPWR VGND sg13g2_decap_4
XFILLER_41_133 VPWR VGND sg13g2_decap_4
X_11661_ _05566_ _05475_ _05434_ VPWR VGND sg13g2_nand2_1
XFILLER_23_870 VPWR VGND sg13g2_fill_1
XFILLER_30_818 VPWR VGND sg13g2_fill_1
X_14380_ _00181_ VGND VPWR _00921_ fpmul.reg_b_out\[11\] clknet_leaf_124_clk sg13g2_dfrbpq_2
X_10612_ _04625_ fp16_res_pipe.add_renorm0.mantisa\[11\] fp16_res_pipe.add_renorm0.mantisa\[6\]
+ VPWR VGND sg13g2_nand2_1
X_11592_ _05491_ _05496_ _05497_ VPWR VGND sg13g2_nor2_1
X_13331_ _07036_ VPWR _00830_ VGND _06980_ net1724 sg13g2_o21ai_1
XFILLER_6_502 VPWR VGND sg13g2_decap_8
X_10543_ _04580_ VPWR _01161_ VGND net1849 _04579_ sg13g2_o21ai_1
XFILLER_10_531 VPWR VGND sg13g2_decap_8
XFILLER_10_542 VPWR VGND sg13g2_fill_1
XFILLER_22_391 VPWR VGND sg13g2_fill_1
XFILLER_127_238 VPWR VGND sg13g2_decap_8
XFILLER_109_942 VPWR VGND sg13g2_decap_8
XFILLER_41_63 VPWR VGND sg13g2_decap_8
XFILLER_108_452 VPWR VGND sg13g2_fill_1
X_13262_ _03272_ _02576_ _06983_ VPWR VGND sg13g2_nor2_1
X_10474_ VGND VPWR _04520_ net1847 _01171_ _04521_ sg13g2_a21oi_1
XFILLER_123_400 VPWR VGND sg13g2_decap_8
X_12213_ _06058_ VPWR _06059_ VGND _06020_ _06057_ sg13g2_o21ai_1
X_13193_ _06930_ net1712 sipo.word\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_6_579 VPWR VGND sg13g2_decap_8
XFILLER_124_956 VPWR VGND sg13g2_decap_8
X_12144_ VPWR _05990_ _05989_ VGND sg13g2_inv_1
XFILLER_111_628 VPWR VGND sg13g2_decap_8
XFILLER_2_752 VPWR VGND sg13g2_fill_1
XFILLER_1_240 VPWR VGND sg13g2_fill_2
XFILLER_104_691 VPWR VGND sg13g2_fill_1
XFILLER_104_680 VPWR VGND sg13g2_decap_8
X_12075_ _05918_ _05920_ _05911_ _05921_ VPWR VGND sg13g2_nand3_1
XFILLER_49_233 VPWR VGND sg13g2_decap_4
XFILLER_2_35 VPWR VGND sg13g2_decap_8
X_11026_ _05003_ _05004_ _05005_ VPWR VGND sg13g2_nor2_1
XFILLER_65_715 VPWR VGND sg13g2_decap_8
XFILLER_38_918 VPWR VGND sg13g2_decap_8
XFILLER_92_578 VPWR VGND sg13g2_decap_8
X_12977_ _06747_ net1717 _00005_ VPWR VGND sg13g2_nand2_1
XFILLER_61_921 VPWR VGND sg13g2_fill_1
XFILLER_61_910 VPWR VGND sg13g2_decap_8
XFILLER_46_984 VPWR VGND sg13g2_fill_1
XFILLER_17_141 VPWR VGND sg13g2_decap_4
XFILLER_18_686 VPWR VGND sg13g2_decap_8
XFILLER_61_954 VPWR VGND sg13g2_decap_8
XFILLER_45_494 VPWR VGND sg13g2_fill_2
X_11928_ _05796_ net1879 fpmul.reg_b_out\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_33_656 VPWR VGND sg13g2_decap_8
X_14716_ _00517_ VGND VPWR _01244_ fp16_res_pipe.exp_mant_logic0.a\[3\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_32_111 VPWR VGND sg13g2_fill_2
XFILLER_33_689 VPWR VGND sg13g2_decap_8
XFILLER_21_818 VPWR VGND sg13g2_fill_2
X_14647_ _00448_ VGND VPWR _01175_ fp16_res_pipe.exp_mant_logic0.b\[0\] clknet_leaf_141_clk
+ sg13g2_dfrbpq_2
X_11859_ VGND VPWR _05754_ _05755_ _05756_ fp16_sum_pipe.seg_reg1.q\[21\] sg13g2_a21oi_1
XFILLER_14_881 VPWR VGND sg13g2_decap_8
X_14578_ _00379_ VGND VPWR _01110_ fp16_sum_pipe.exp_mant_logic0.b\[5\] clknet_leaf_117_clk
+ sg13g2_dfrbpq_1
X_13529_ VPWR _00080_ net84 VGND sg13g2_inv_1
XFILLER_118_238 VPWR VGND sg13g2_decap_8
XFILLER_9_373 VPWR VGND sg13g2_decap_8
XFILLER_127_750 VPWR VGND sg13g2_decap_8
XFILLER_115_956 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_114_466 VPWR VGND sg13g2_fill_2
XFILLER_114_455 VPWR VGND sg13g2_decap_8
X_07952_ VPWR _02226_ fp16_sum_pipe.seg_reg0.q\[28\] VGND sg13g2_inv_1
X_07883_ _02168_ VPWR _01402_ VGND net1895 _01825_ sg13g2_o21ai_1
XFILLER_96_873 VPWR VGND sg13g2_decap_8
XFILLER_68_575 VPWR VGND sg13g2_decap_8
XFILLER_68_564 VPWR VGND sg13g2_fill_1
X_09622_ _03737_ _03738_ _03736_ _03739_ VPWR VGND sg13g2_nand3_1
XFILLER_83_534 VPWR VGND sg13g2_fill_1
XFILLER_83_523 VPWR VGND sg13g2_decap_8
XFILLER_83_512 VPWR VGND sg13g2_fill_1
XFILLER_56_748 VPWR VGND sg13g2_decap_8
XFILLER_56_737 VPWR VGND sg13g2_fill_2
X_09553_ VPWR _03670_ acc_sum.add_renorm0.mantisa\[2\] VGND sg13g2_inv_1
XFILLER_83_545 VPWR VGND sg13g2_fill_2
XFILLER_55_236 VPWR VGND sg13g2_fill_2
XFILLER_102_14 VPWR VGND sg13g2_decap_8
X_08504_ VGND VPWR net1740 net1816 _01348_ _02728_ sg13g2_a21oi_1
XFILLER_37_973 VPWR VGND sg13g2_decap_8
XFILLER_36_494 VPWR VGND sg13g2_decap_8
X_09484_ _03607_ net1828 VPWR VGND sg13g2_inv_2
X_08435_ _02669_ fpdiv.divider0.divisor_reg\[7\] fpdiv.divider0.remainder_reg\[7\]
+ VPWR VGND sg13g2_xnor2_1
XFILLER_52_987 VPWR VGND sg13g2_decap_8
XFILLER_23_133 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_fill_2
X_08366_ _02606_ instr\[2\] _02608_ _02609_ VPWR VGND sg13g2_nor3_1
XFILLER_51_497 VPWR VGND sg13g2_decap_8
XFILLER_23_188 VPWR VGND sg13g2_fill_2
XFILLER_23_199 VPWR VGND sg13g2_decap_8
X_07317_ _01681_ net1784 acc_sub.add_renorm0.mantisa\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_20_840 VPWR VGND sg13g2_decap_8
XFILLER_127_7 VPWR VGND sg13g2_decap_8
X_08297_ _02541_ _02542_ _02543_ _02544_ VPWR VGND sg13g2_nor3_1
X_07248_ _01619_ net1784 acc_sub.add_renorm0.mantisa\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_118_761 VPWR VGND sg13g2_decap_8
XFILLER_109_249 VPWR VGND sg13g2_decap_4
XFILLER_106_901 VPWR VGND sg13g2_decap_8
X_07179_ _01551_ _01550_ acc_sub.op_sign_logic0.mantisa_a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_106_978 VPWR VGND sg13g2_decap_8
XFILLER_105_422 VPWR VGND sg13g2_fill_1
XFILLER_11_77 VPWR VGND sg13g2_decap_8
X_10190_ _04265_ _04266_ _04264_ _04268_ VPWR VGND _04267_ sg13g2_nand4_1
XFILLER_127_77 VPWR VGND sg13g2_decap_8
XFILLER_121_959 VPWR VGND sg13g2_decap_8
XFILLER_120_447 VPWR VGND sg13g2_decap_4
XFILLER_105_499 VPWR VGND sg13g2_decap_8
XFILLER_87_862 VPWR VGND sg13g2_fill_1
XFILLER_87_851 VPWR VGND sg13g2_fill_2
XFILLER_86_350 VPWR VGND sg13g2_decap_8
XFILLER_59_553 VPWR VGND sg13g2_fill_1
XFILLER_59_542 VPWR VGND sg13g2_decap_8
XFILLER_4_1007 VPWR VGND sg13g2_decap_8
XFILLER_101_694 VPWR VGND sg13g2_fill_1
XFILLER_74_512 VPWR VGND sg13g2_decap_8
X_12900_ _06676_ _06672_ _06675_ _06510_ net1948 VPWR VGND sg13g2_a22oi_1
X_13880_ VPWR _00431_ net48 VGND sg13g2_inv_1
X_12831_ _06613_ _06612_ net1732 VPWR VGND sg13g2_nand2_1
XFILLER_46_225 VPWR VGND sg13g2_decap_8
XFILLER_62_729 VPWR VGND sg13g2_decap_8
XFILLER_43_921 VPWR VGND sg13g2_decap_4
XFILLER_36_63 VPWR VGND sg13g2_decap_8
XFILLER_28_973 VPWR VGND sg13g2_decap_8
X_12762_ _06547_ net1767 acc\[15\] net1908 VPWR VGND sg13g2_and3_1
X_14501_ _00302_ VGND VPWR _01037_ fpdiv.reg_b_out\[8\] clknet_leaf_54_clk sg13g2_dfrbpq_1
X_12693_ VPWR _06502_ div_result\[7\] VGND sg13g2_inv_1
XFILLER_70_773 VPWR VGND sg13g2_decap_8
XFILLER_15_667 VPWR VGND sg13g2_decap_8
X_11713_ _05617_ _05616_ VPWR VGND sg13g2_inv_2
X_14432_ _00233_ VGND VPWR _00971_ fpmul.seg_reg0.q\[17\] clknet_leaf_101_clk sg13g2_dfrbpq_1
XFILLER_42_497 VPWR VGND sg13g2_fill_2
X_11644_ _05549_ _05548_ _05498_ VPWR VGND sg13g2_nand2_1
XFILLER_122_1012 VPWR VGND sg13g2_fill_2
XFILLER_122_1001 VPWR VGND sg13g2_decap_8
XFILLER_11_840 VPWR VGND sg13g2_decap_8
X_14363_ _00164_ VGND VPWR _00905_ _00016_ clknet_leaf_87_clk sg13g2_dfrbpq_1
X_11575_ net1836 VPWR _05480_ VGND _05463_ _05479_ sg13g2_o21ai_1
X_14294_ _00095_ VGND VPWR _00838_ acc\[4\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_13314_ _07024_ net1742 sipo.word\[0\] VPWR VGND sg13g2_nand2_1
X_10526_ _04567_ _04428_ _04566_ VPWR VGND sg13g2_xnor2_1
X_13245_ _06969_ VPWR _00849_ VGND _01723_ _06962_ sg13g2_o21ai_1
XFILLER_7_888 VPWR VGND sg13g2_decap_8
X_10457_ _04505_ _04504_ _04458_ VPWR VGND sg13g2_nand2_1
XFILLER_124_753 VPWR VGND sg13g2_decap_8
XFILLER_6_398 VPWR VGND sg13g2_decap_4
XFILLER_123_252 VPWR VGND sg13g2_decap_8
XFILLER_112_915 VPWR VGND sg13g2_decap_8
XFILLER_97_626 VPWR VGND sg13g2_fill_1
XFILLER_69_317 VPWR VGND sg13g2_decap_8
X_13176_ VPWR _06918_ sipo.shift_reg\[12\] VGND sg13g2_inv_1
XFILLER_42_7 VPWR VGND sg13g2_decap_8
X_10388_ VPWR _04438_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[5\] VGND sg13g2_inv_1
XFILLER_111_436 VPWR VGND sg13g2_decap_8
XFILLER_78_840 VPWR VGND sg13g2_decap_8
X_12127_ VGND VPWR _05965_ _05971_ _05973_ _05972_ sg13g2_a21oi_1
XFILLER_111_447 VPWR VGND sg13g2_fill_1
XFILLER_84_309 VPWR VGND sg13g2_decap_8
XFILLER_78_873 VPWR VGND sg13g2_decap_4
X_12058_ _05903_ VPWR _05904_ VGND _05899_ _05900_ sg13g2_o21ai_1
XFILLER_42_1013 VPWR VGND sg13g2_fill_1
XFILLER_38_704 VPWR VGND sg13g2_decap_8
XFILLER_120_981 VPWR VGND sg13g2_decap_8
XFILLER_77_361 VPWR VGND sg13g2_fill_2
XFILLER_38_726 VPWR VGND sg13g2_fill_1
XFILLER_37_214 VPWR VGND sg13g2_fill_2
X_11009_ _04990_ VPWR _01105_ VGND net1929 _02469_ sg13g2_o21ai_1
XFILLER_93_854 VPWR VGND sg13g2_decap_8
XFILLER_65_534 VPWR VGND sg13g2_decap_8
XFILLER_37_225 VPWR VGND sg13g2_decap_8
XFILLER_93_898 VPWR VGND sg13g2_decap_8
XFILLER_92_353 VPWR VGND sg13g2_decap_8
XFILLER_53_729 VPWR VGND sg13g2_fill_2
XFILLER_80_559 VPWR VGND sg13g2_fill_1
XFILLER_34_954 VPWR VGND sg13g2_decap_8
X_08220_ _02351_ _02250_ _02475_ VPWR VGND sg13g2_nor2b_1
XFILLER_33_497 VPWR VGND sg13g2_fill_2
X_08151_ _02410_ VPWR _02411_ VGND _02268_ net1648 sg13g2_o21ai_1
XFILLER_119_558 VPWR VGND sg13g2_decap_8
XFILLER_107_709 VPWR VGND sg13g2_fill_1
XFILLER_106_208 VPWR VGND sg13g2_fill_2
XFILLER_115_753 VPWR VGND sg13g2_decap_8
XFILLER_114_263 VPWR VGND sg13g2_decap_8
XFILLER_0_519 VPWR VGND sg13g2_decap_8
X_08984_ _03169_ _03139_ _03170_ VPWR VGND sg13g2_and2_1
XFILLER_88_637 VPWR VGND sg13g2_decap_8
XFILLER_57_18 VPWR VGND sg13g2_fill_1
X_07935_ _02210_ fp16_sum_pipe.exp_mant_logic0.b\[9\] VPWR VGND sg13g2_inv_2
XFILLER_111_992 VPWR VGND sg13g2_decap_8
XFILLER_96_692 VPWR VGND sg13g2_decap_4
XFILLER_28_214 VPWR VGND sg13g2_decap_8
XFILLER_113_35 VPWR VGND sg13g2_decap_8
X_09605_ VGND VPWR _03689_ net1804 _03722_ _03721_ sg13g2_a21oi_1
X_07866_ _02160_ _02159_ _02063_ VPWR VGND sg13g2_nand2_1
XFILLER_84_865 VPWR VGND sg13g2_fill_2
XFILLER_83_342 VPWR VGND sg13g2_fill_1
XFILLER_68_394 VPWR VGND sg13g2_fill_2
X_07797_ VPWR _02096_ acc_sub.exp_mant_logic0.b\[6\] VGND sg13g2_inv_1
XFILLER_83_375 VPWR VGND sg13g2_fill_1
XFILLER_71_504 VPWR VGND sg13g2_fill_1
XFILLER_56_567 VPWR VGND sg13g2_decap_8
XFILLER_37_770 VPWR VGND sg13g2_fill_2
XFILLER_16_409 VPWR VGND sg13g2_fill_1
XFILLER_25_910 VPWR VGND sg13g2_decap_8
XFILLER_83_397 VPWR VGND sg13g2_decap_8
XFILLER_71_559 VPWR VGND sg13g2_decap_8
XFILLER_43_228 VPWR VGND sg13g2_decap_8
X_09467_ _03596_ acc_sub.x2\[11\] net1914 VPWR VGND sg13g2_nand2_1
XFILLER_36_291 VPWR VGND sg13g2_decap_4
XFILLER_25_987 VPWR VGND sg13g2_decap_8
XFILLER_51_250 VPWR VGND sg13g2_fill_1
XFILLER_40_924 VPWR VGND sg13g2_decap_8
X_09398_ VGND VPWR _03543_ _03425_ _03544_ _03518_ sg13g2_a21oi_1
X_08349_ _02592_ _02591_ VPWR VGND sg13g2_inv_2
XFILLER_22_21 VPWR VGND sg13g2_decap_8
X_11360_ _05311_ VPWR _05312_ VGND _03353_ _05143_ sg13g2_o21ai_1
X_10311_ _04373_ net1912 fp16_res_pipe.x2\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_4_825 VPWR VGND sg13g2_decap_8
X_13030_ VGND VPWR _06750_ fpmul.seg_reg0.q\[4\] _06798_ fpmul.seg_reg0.q\[5\] sg13g2_a21oi_1
X_11291_ _03351_ _03353_ _03345_ _05251_ VPWR VGND _03357_ sg13g2_nand4_1
XFILLER_3_335 VPWR VGND sg13g2_decap_4
XFILLER_3_324 VPWR VGND sg13g2_decap_8
XFILLER_121_701 VPWR VGND sg13g2_fill_1
XFILLER_105_241 VPWR VGND sg13g2_decap_4
X_10242_ _04314_ net1688 fp16_res_pipe.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
X_10173_ _04253_ _04252_ net1637 VPWR VGND sg13g2_nand2_1
XFILLER_121_756 VPWR VGND sg13g2_decap_8
XFILLER_78_147 VPWR VGND sg13g2_decap_8
XFILLER_120_266 VPWR VGND sg13g2_decap_8
XFILLER_93_117 VPWR VGND sg13g2_decap_8
XFILLER_87_670 VPWR VGND sg13g2_fill_2
XFILLER_47_501 VPWR VGND sg13g2_fill_1
XFILLER_47_40 VPWR VGND sg13g2_decap_8
XFILLER_47_545 VPWR VGND sg13g2_decap_8
X_13932_ VPWR _00483_ net5 VGND sg13g2_inv_1
XFILLER_35_707 VPWR VGND sg13g2_decap_8
X_13863_ VPWR _00414_ net51 VGND sg13g2_inv_1
XFILLER_16_910 VPWR VGND sg13g2_decap_8
XFILLER_90_846 VPWR VGND sg13g2_decap_4
X_12814_ _06596_ _06595_ net1923 _06597_ VPWR VGND sg13g2_a21o_1
X_13794_ VPWR _00345_ net20 VGND sg13g2_inv_1
XFILLER_28_792 VPWR VGND sg13g2_decap_8
Xclkbuf_5_21__f_clk clknet_4_10_0_clk clknet_5_21__leaf_clk VPWR VGND sg13g2_buf_8
X_12745_ fpmul.reg_b_out\[12\] fp16_res_pipe.x2\[12\] net1952 _00922_ VPWR VGND sg13g2_mux2_1
XFILLER_15_431 VPWR VGND sg13g2_fill_1
XFILLER_16_987 VPWR VGND sg13g2_decap_8
XFILLER_43_773 VPWR VGND sg13g2_fill_1
XFILLER_42_261 VPWR VGND sg13g2_fill_2
XFILLER_31_935 VPWR VGND sg13g2_decap_8
X_12676_ _06354_ net1735 _06489_ VPWR VGND sg13g2_nor2_1
XFILLER_30_445 VPWR VGND sg13g2_fill_1
X_14415_ _00216_ VGND VPWR _00954_ fpmul.reg_a_out\[12\] clknet_leaf_127_clk sg13g2_dfrbpq_2
XFILLER_8_56 VPWR VGND sg13g2_decap_8
X_11627_ _05532_ _05526_ _05531_ VPWR VGND sg13g2_xnor2_1
X_14346_ _00147_ VGND VPWR _00888_ fpmul.reg_p_out\[10\] clknet_leaf_88_clk sg13g2_dfrbpq_1
X_11558_ _05430_ _05435_ _05462_ _05463_ VPWR VGND sg13g2_nor3_1
XFILLER_116_528 VPWR VGND sg13g2_decap_8
XFILLER_7_685 VPWR VGND sg13g2_decap_8
XFILLER_6_140 VPWR VGND sg13g2_decap_8
X_10509_ _04552_ net1673 _04551_ VPWR VGND sg13g2_nand2b_1
X_11489_ _05397_ VPWR _01032_ VGND net1945 _01768_ sg13g2_o21ai_1
X_14277_ _00078_ VGND VPWR _00828_ fp16_res_pipe.x2\[10\] clknet_leaf_128_clk sg13g2_dfrbpq_2
XFILLER_7_696 VPWR VGND sg13g2_fill_2
X_13228_ sipo.word_ready _06952_ _06953_ VPWR VGND sg13g2_nor2_1
XFILLER_98_946 VPWR VGND sg13g2_decap_8
XFILLER_88_91 VPWR VGND sg13g2_decap_8
XFILLER_69_114 VPWR VGND sg13g2_fill_2
X_13159_ _06905_ _06903_ VPWR VGND sg13g2_inv_2
XFILLER_97_456 VPWR VGND sg13g2_fill_2
XFILLER_112_789 VPWR VGND sg13g2_decap_8
XFILLER_111_288 VPWR VGND sg13g2_decap_8
XFILLER_111_277 VPWR VGND sg13g2_fill_2
X_07720_ _02023_ _02026_ _02027_ VPWR VGND sg13g2_nor2_1
XFILLER_97_478 VPWR VGND sg13g2_decap_4
XFILLER_66_843 VPWR VGND sg13g2_fill_2
XFILLER_65_331 VPWR VGND sg13g2_fill_2
X_07651_ _01963_ _01958_ _01962_ VPWR VGND sg13g2_nand2_1
XFILLER_80_301 VPWR VGND sg13g2_decap_8
XFILLER_65_353 VPWR VGND sg13g2_decap_8
XFILLER_53_504 VPWR VGND sg13g2_fill_1
XFILLER_92_161 VPWR VGND sg13g2_decap_8
X_07582_ _01896_ _01787_ _01895_ VPWR VGND sg13g2_xnor2_1
XFILLER_53_526 VPWR VGND sg13g2_decap_8
XFILLER_19_792 VPWR VGND sg13g2_decap_8
X_09321_ _03473_ VPWR _03474_ VGND _03378_ _03380_ sg13g2_o21ai_1
XFILLER_80_389 VPWR VGND sg13g2_fill_2
XFILLER_61_570 VPWR VGND sg13g2_decap_4
XFILLER_34_784 VPWR VGND sg13g2_decap_4
XFILLER_33_250 VPWR VGND sg13g2_decap_8
X_09252_ fp16_res_pipe.op_sign_logic0.mantisa_b\[2\] _03405_ _03406_ VPWR VGND sg13g2_nor2_1
XFILLER_22_968 VPWR VGND sg13g2_decap_8
X_09183_ _03345_ acc_sum.exp_mant_logic0.b\[6\] VPWR VGND sg13g2_inv_2
X_08203_ _02459_ fp16_sum_pipe.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_inv_2
XFILLER_88_1013 VPWR VGND sg13g2_fill_1
XFILLER_88_1002 VPWR VGND sg13g2_decap_8
X_08134_ _02392_ _02393_ _02394_ _02395_ VPWR VGND sg13g2_nor3_1
XFILLER_30_990 VPWR VGND sg13g2_decap_8
XFILLER_119_377 VPWR VGND sg13g2_decap_8
XFILLER_108_35 VPWR VGND sg13g2_fill_2
Xplace1830 fp16_res_pipe.exp_mant_logic0.b\[5\] net1830 VPWR VGND sg13g2_buf_2
X_08065_ _02221_ _02326_ _02311_ _02331_ VPWR VGND sg13g2_nor3_1
XFILLER_122_509 VPWR VGND sg13g2_fill_1
Xplace1852 net1851 net1852 VPWR VGND sg13g2_buf_2
Xplace1863 fpmul.reg_b_out\[6\] net1863 VPWR VGND sg13g2_buf_2
Xplace1841 fp16_sum_pipe.add_renorm0.mantisa\[11\] net1841 VPWR VGND sg13g2_buf_1
XFILLER_88_434 VPWR VGND sg13g2_decap_8
Xplace1885 acc_sub.reg1en.d\[0\] net1885 VPWR VGND sg13g2_buf_2
Xplace1896 acc_sum.reg1en.d\[0\] net1896 VPWR VGND sg13g2_buf_2
Xplace1874 net1873 net1874 VPWR VGND sg13g2_buf_2
XFILLER_102_233 VPWR VGND sg13g2_decap_8
XFILLER_102_222 VPWR VGND sg13g2_decap_4
XFILLER_89_979 VPWR VGND sg13g2_decap_8
XFILLER_88_456 VPWR VGND sg13g2_decap_8
XFILLER_76_607 VPWR VGND sg13g2_fill_2
XFILLER_124_56 VPWR VGND sg13g2_decap_8
X_08967_ VGND VPWR _03152_ _03153_ _03151_ net1699 sg13g2_a21oi_2
XFILLER_76_618 VPWR VGND sg13g2_decap_8
XFILLER_57_821 VPWR VGND sg13g2_decap_8
XFILLER_48_309 VPWR VGND sg13g2_fill_2
XFILLER_29_501 VPWR VGND sg13g2_fill_2
X_08898_ _02991_ _02998_ _03085_ VPWR VGND sg13g2_nor2_1
XFILLER_57_832 VPWR VGND sg13g2_fill_1
X_07918_ fp16_sum_pipe.exp_mant_logic0.b\[11\] _02192_ _02193_ VPWR VGND sg13g2_nor2_1
X_07849_ _02144_ _02142_ _02143_ VPWR VGND sg13g2_nand2_1
XFILLER_72_813 VPWR VGND sg13g2_decap_8
XFILLER_56_364 VPWR VGND sg13g2_fill_2
XFILLER_17_21 VPWR VGND sg13g2_decap_8
X_10860_ net1824 fp16_res_pipe.add_renorm0.exp\[3\] _04872_ VPWR VGND sg13g2_nor2_1
XFILLER_71_356 VPWR VGND sg13g2_decap_8
XFILLER_24_261 VPWR VGND sg13g2_decap_8
XFILLER_24_272 VPWR VGND sg13g2_fill_1
X_10791_ VPWR _04803_ fp16_res_pipe.add_renorm0.exp\[0\] VGND sg13g2_inv_1
X_12530_ _06351_ acc_sub.x2\[2\] net1954 VPWR VGND sg13g2_nand2_1
XFILLER_9_906 VPWR VGND sg13g2_decap_8
XFILLER_12_434 VPWR VGND sg13g2_fill_2
XFILLER_13_968 VPWR VGND sg13g2_decap_8
XFILLER_33_42 VPWR VGND sg13g2_decap_8
X_12461_ _06303_ VPWR _00966_ VGND net1870 _06301_ sg13g2_o21ai_1
XFILLER_33_86 VPWR VGND sg13g2_fill_1
X_14200_ VPWR _00751_ net105 VGND sg13g2_inv_1
X_11412_ _05352_ net1718 fpdiv.div_out\[1\] VPWR VGND sg13g2_nand2_1
X_14131_ VPWR _00682_ net103 VGND sg13g2_inv_1
X_12392_ VPWR _06238_ _06237_ VGND sg13g2_inv_1
XFILLER_126_848 VPWR VGND sg13g2_decap_8
X_11343_ _01077_ _05295_ _05296_ VPWR VGND sg13g2_nand2_1
X_14062_ VPWR _00613_ net94 VGND sg13g2_inv_1
X_11274_ _05234_ _05235_ _05233_ _05236_ VPWR VGND sg13g2_nand3_1
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_106_572 VPWR VGND sg13g2_fill_2
X_13013_ _06777_ _06779_ _06781_ VPWR VGND sg13g2_nor2_1
X_10225_ fp16_res_pipe.exp_mant_logic0.b\[2\] _04298_ VPWR VGND sg13g2_inv_4
XFILLER_66_117 VPWR VGND sg13g2_decap_8
X_10156_ _04237_ net1643 fp16_res_pipe.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
X_14964_ _00765_ VGND VPWR _01484_ acc_sub.add_renorm0.mantisa\[8\] clknet_leaf_63_clk
+ sg13g2_dfrbpq_2
XFILLER_75_640 VPWR VGND sg13g2_decap_8
XFILLER_48_843 VPWR VGND sg13g2_fill_1
X_10087_ VGND VPWR fp16_res_pipe.exp_mant_logic0.a\[4\] _04126_ _04172_ _04171_ sg13g2_a21oi_1
XFILLER_35_504 VPWR VGND sg13g2_decap_8
X_13915_ VPWR _00466_ net5 VGND sg13g2_inv_1
X_14895_ _00696_ VGND VPWR _01415_ acc_sub.op_sign_logic0.mantisa_b\[5\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_1
XFILLER_74_60 VPWR VGND sg13g2_decap_8
XFILLER_90_654 VPWR VGND sg13g2_decap_8
XFILLER_63_868 VPWR VGND sg13g2_decap_8
X_13846_ VPWR _00397_ net29 VGND sg13g2_inv_1
X_13777_ VPWR _00328_ net139 VGND sg13g2_inv_1
X_10989_ _04980_ VPWR _01115_ VGND net1931 _02205_ sg13g2_o21ai_1
X_12728_ _06532_ VPWR _00929_ VGND _06527_ _02648_ sg13g2_o21ai_1
XFILLER_43_581 VPWR VGND sg13g2_decap_8
X_12659_ _06475_ _06472_ _06474_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_798 VPWR VGND sg13g2_decap_8
XFILLER_117_837 VPWR VGND sg13g2_decap_8
XFILLER_8_972 VPWR VGND sg13g2_decap_8
X_14329_ _00130_ VGND VPWR _00003_ sipo.receiving clknet_leaf_8_clk sg13g2_dfrbpq_1
X_09870_ _03976_ _03649_ _03652_ VPWR VGND sg13g2_nand2_1
X_08821_ _03008_ _03001_ _03007_ _02999_ _02967_ VPWR VGND sg13g2_a22oi_1
XFILLER_97_220 VPWR VGND sg13g2_fill_2
XFILLER_31_0 VPWR VGND sg13g2_decap_8
XFILLER_97_286 VPWR VGND sg13g2_decap_4
XFILLER_86_938 VPWR VGND sg13g2_decap_8
XFILLER_100_737 VPWR VGND sg13g2_decap_8
X_08752_ _02948_ acc\[8\] net1900 VPWR VGND sg13g2_nand2_1
XFILLER_39_854 VPWR VGND sg13g2_decap_8
XFILLER_38_331 VPWR VGND sg13g2_decap_4
X_07703_ _02011_ _02004_ _02010_ VPWR VGND sg13g2_nand2_1
XFILLER_94_982 VPWR VGND sg13g2_decap_8
X_08683_ _02899_ _02774_ _02898_ VPWR VGND sg13g2_xnor2_1
X_07634_ _01948_ net1792 net1672 acc_sub.op_sign_logic0.mantisa_a\[9\] net1779 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_93_481 VPWR VGND sg13g2_decap_4
XFILLER_66_695 VPWR VGND sg13g2_decap_8
XFILLER_65_172 VPWR VGND sg13g2_fill_2
XFILLER_65_161 VPWR VGND sg13g2_fill_1
XFILLER_53_312 VPWR VGND sg13g2_fill_2
XFILLER_0_1010 VPWR VGND sg13g2_decap_4
XFILLER_81_643 VPWR VGND sg13g2_fill_1
XFILLER_54_879 VPWR VGND sg13g2_fill_1
XFILLER_26_559 VPWR VGND sg13g2_decap_8
XFILLER_110_14 VPWR VGND sg13g2_decap_8
X_07565_ _01879_ _01878_ _01790_ VPWR VGND sg13g2_nand2b_1
XFILLER_55_1012 VPWR VGND sg13g2_fill_2
X_07496_ VPWR _01819_ _01818_ VGND sg13g2_inv_1
X_09304_ _03457_ VPWR _03458_ VGND fp16_res_pipe.op_sign_logic0.s_a _03453_ sg13g2_o21ai_1
XFILLER_22_732 VPWR VGND sg13g2_decap_4
XFILLER_22_743 VPWR VGND sg13g2_fill_2
X_09235_ VPWR _03389_ _03388_ VGND sg13g2_inv_1
XFILLER_10_905 VPWR VGND sg13g2_decap_8
XFILLER_22_787 VPWR VGND sg13g2_fill_1
XFILLER_108_826 VPWR VGND sg13g2_fill_1
X_09166_ _03334_ acc_sub.x2\[12\] net1904 VPWR VGND sg13g2_nand2_1
XFILLER_119_196 VPWR VGND sg13g2_decap_8
XFILLER_119_56 VPWR VGND sg13g2_decap_8
X_09097_ _03280_ _03233_ _03231_ VPWR VGND sg13g2_xnor2_1
X_08048_ _02313_ _02212_ _02314_ VPWR VGND sg13g2_xor2_1
XFILLER_116_870 VPWR VGND sg13g2_decap_8
Xplace1660 _01905_ net1660 VPWR VGND sg13g2_buf_2
XFILLER_89_732 VPWR VGND sg13g2_decap_8
Xplace1671 _02800_ net1671 VPWR VGND sg13g2_buf_2
XFILLER_103_542 VPWR VGND sg13g2_decap_8
Xplace1693 _07055_ net1693 VPWR VGND sg13g2_buf_2
XFILLER_49_607 VPWR VGND sg13g2_decap_8
X_10010_ _04098_ _04050_ _04086_ VPWR VGND sg13g2_nand2_1
Xplace1682 _04056_ net1682 VPWR VGND sg13g2_buf_2
XFILLER_89_787 VPWR VGND sg13g2_decap_8
XFILLER_88_275 VPWR VGND sg13g2_fill_1
XFILLER_77_927 VPWR VGND sg13g2_decap_4
XFILLER_49_618 VPWR VGND sg13g2_fill_2
X_09999_ VGND VPWR _04086_ _04042_ _04087_ _03996_ sg13g2_a21oi_1
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_88_297 VPWR VGND sg13g2_fill_2
XFILLER_88_286 VPWR VGND sg13g2_decap_8
XFILLER_85_971 VPWR VGND sg13g2_decap_8
XFILLER_63_109 VPWR VGND sg13g2_decap_4
X_11961_ _05818_ net1884 fpmul.reg_b_out\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_28_42 VPWR VGND sg13g2_decap_8
XFILLER_72_632 VPWR VGND sg13g2_fill_2
X_13700_ VPWR _00251_ net54 VGND sg13g2_inv_1
X_10912_ _04915_ _04888_ _04921_ VPWR VGND sg13g2_nor2_1
XFILLER_72_654 VPWR VGND sg13g2_decap_8
XFILLER_71_120 VPWR VGND sg13g2_decap_8
XFILLER_60_805 VPWR VGND sg13g2_fill_1
X_11892_ _05777_ fpmul.reg_a_out\[15\] fpmul.reg_b_out\[15\] VPWR VGND sg13g2_xnor2_1
X_14680_ _00481_ VGND VPWR _01208_ fp16_res_pipe.op_sign_logic0.mantisa_a\[6\] clknet_leaf_144_clk
+ sg13g2_dfrbpq_2
X_13631_ VPWR _00182_ net50 VGND sg13g2_inv_1
X_10843_ _04854_ _04737_ _04853_ _04855_ VPWR VGND sg13g2_nand3_1
X_13562_ VPWR _00113_ net83 VGND sg13g2_inv_1
XFILLER_44_63 VPWR VGND sg13g2_decap_8
X_10774_ fp16_res_pipe.add_renorm0.mantisa\[10\] fp16_res_pipe.add_renorm0.mantisa\[9\]
+ _04651_ _04786_ VPWR VGND sg13g2_nand3_1
XFILLER_12_220 VPWR VGND sg13g2_fill_1
X_12513_ fpmul.reg_a_out\[10\] net1953 _06342_ VPWR VGND sg13g2_nor2_1
XFILLER_9_736 VPWR VGND sg13g2_fill_1
X_13493_ VPWR _00044_ net32 VGND sg13g2_inv_1
XFILLER_40_584 VPWR VGND sg13g2_decap_8
XFILLER_12_286 VPWR VGND sg13g2_decap_4
X_12444_ _06290_ _06287_ _06286_ VPWR VGND sg13g2_nand2b_1
XFILLER_60_62 VPWR VGND sg13g2_fill_2
XFILLER_60_51 VPWR VGND sg13g2_fill_2
X_12375_ _06221_ _06217_ _06218_ VPWR VGND sg13g2_xnor2_1
XFILLER_60_95 VPWR VGND sg13g2_decap_4
XFILLER_5_920 VPWR VGND sg13g2_decap_8
XFILLER_125_133 VPWR VGND sg13g2_decap_8
XFILLER_114_818 VPWR VGND sg13g2_decap_8
X_11326_ _05252_ _05183_ _05281_ VPWR VGND sg13g2_nor2_1
X_14114_ VPWR _00665_ net44 VGND sg13g2_inv_1
XFILLER_5_35 VPWR VGND sg13g2_decap_8
XFILLER_4_441 VPWR VGND sg13g2_decap_8
X_14045_ VPWR _00596_ net76 VGND sg13g2_inv_1
XFILLER_5_997 VPWR VGND sg13g2_decap_8
XFILLER_122_840 VPWR VGND sg13g2_decap_8
X_11257_ _05220_ net1661 acc_sum.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_69_82 VPWR VGND sg13g2_fill_1
X_11188_ _05155_ _05156_ _05154_ _05157_ VPWR VGND sg13g2_nand3_1
XFILLER_68_938 VPWR VGND sg13g2_decap_8
XFILLER_67_404 VPWR VGND sg13g2_fill_2
X_10208_ _04283_ _04165_ net1745 VPWR VGND sg13g2_nand2_1
XFILLER_79_286 VPWR VGND sg13g2_fill_2
XFILLER_0_691 VPWR VGND sg13g2_decap_8
X_10139_ _04221_ fp16_res_pipe.exp_mant_logic0.a\[0\] net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[3\]
+ net1763 VPWR VGND sg13g2_a22oi_1
XFILLER_94_256 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_fill_1
XFILLER_36_802 VPWR VGND sg13g2_decap_8
X_14947_ _00748_ VGND VPWR _01467_ acc_sub.exp_mant_logic0.a\[15\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_2
XFILLER_85_92 VPWR VGND sg13g2_fill_1
XFILLER_75_481 VPWR VGND sg13g2_fill_2
XFILLER_75_470 VPWR VGND sg13g2_decap_4
X_14878_ _00679_ VGND VPWR _01398_ acc_sub.exp_mant_logic0.b\[4\] clknet_leaf_58_clk
+ sg13g2_dfrbpq_2
XFILLER_51_805 VPWR VGND sg13g2_decap_8
XFILLER_36_879 VPWR VGND sg13g2_fill_2
XFILLER_36_868 VPWR VGND sg13g2_fill_2
XFILLER_91_996 VPWR VGND sg13g2_decap_8
XFILLER_90_484 VPWR VGND sg13g2_fill_2
XFILLER_63_687 VPWR VGND sg13g2_decap_4
X_13829_ VPWR _00380_ net10 VGND sg13g2_inv_1
X_07350_ VPWR _01709_ acc_sub.add_renorm0.exp\[7\] VGND sg13g2_inv_1
XFILLER_31_562 VPWR VGND sg13g2_decap_8
X_09020_ VPWR _03206_ _03157_ VGND sg13g2_inv_1
X_07281_ VPWR _01649_ _01612_ VGND sg13g2_inv_1
XFILLER_79_0 VPWR VGND sg13g2_decap_4
XFILLER_117_623 VPWR VGND sg13g2_decap_8
XFILLER_116_166 VPWR VGND sg13g2_decap_8
XFILLER_105_829 VPWR VGND sg13g2_decap_8
XFILLER_113_851 VPWR VGND sg13g2_decap_8
XFILLER_59_905 VPWR VGND sg13g2_fill_1
X_09922_ _04019_ _04018_ fp16_res_pipe.exp_mant_logic0.a\[10\] VPWR VGND sg13g2_nand2_1
X_09853_ net1664 _03962_ _03963_ VPWR VGND _03847_ sg13g2_nand3b_1
X_08804_ _02991_ net1704 _02990_ VPWR VGND sg13g2_nand2_1
XFILLER_112_372 VPWR VGND sg13g2_fill_1
XFILLER_100_512 VPWR VGND sg13g2_fill_2
X_09784_ net1769 VPWR _03899_ VGND _03897_ _03898_ sg13g2_o21ai_1
XFILLER_58_448 VPWR VGND sg13g2_decap_4
XFILLER_73_407 VPWR VGND sg13g2_fill_1
X_08735_ _02936_ VPWR _01325_ VGND net1903 _02935_ sg13g2_o21ai_1
XFILLER_27_846 VPWR VGND sg13g2_decap_8
XFILLER_121_35 VPWR VGND sg13g2_decap_8
X_08666_ VGND VPWR net1671 _02876_ _02884_ net1740 sg13g2_a21oi_1
XFILLER_81_440 VPWR VGND sg13g2_fill_2
XFILLER_66_492 VPWR VGND sg13g2_decap_8
X_07617_ VGND VPWR _01927_ _01929_ _01931_ net1660 sg13g2_a21oi_1
XFILLER_92_1009 VPWR VGND sg13g2_decap_4
XFILLER_82_996 VPWR VGND sg13g2_decap_8
X_08597_ VPWR _02820_ _02819_ VGND sg13g2_inv_1
XFILLER_42_838 VPWR VGND sg13g2_fill_2
XFILLER_26_367 VPWR VGND sg13g2_decap_8
X_07548_ _01863_ VPWR _01432_ VGND _01813_ _01855_ sg13g2_o21ai_1
XFILLER_35_890 VPWR VGND sg13g2_decap_8
XFILLER_22_562 VPWR VGND sg13g2_decap_4
X_07479_ _01802_ _01793_ _01797_ _01801_ VPWR VGND sg13g2_and3_1
XFILLER_14_77 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_142_clk clknet_5_0__leaf_clk clknet_leaf_142_clk VPWR VGND sg13g2_buf_8
X_10490_ VGND VPWR _04534_ net1847 _01169_ _04535_ sg13g2_a21oi_1
X_09218_ VPWR _03372_ fp16_res_pipe.op_sign_logic0.mantisa_a\[9\] VGND sg13g2_inv_1
X_09149_ VGND VPWR _03120_ acc_sub.reg3en.q\[0\] _01298_ _03323_ sg13g2_a21oi_1
XFILLER_30_21 VPWR VGND sg13g2_decap_8
XFILLER_107_133 VPWR VGND sg13g2_decap_8
X_12160_ _06006_ _06003_ _06004_ VPWR VGND sg13g2_nand2_1
XFILLER_108_689 VPWR VGND sg13g2_decap_8
X_11111_ VGND VPWR _05033_ _05016_ _05081_ _05013_ sg13g2_a21oi_1
XFILLER_2_912 VPWR VGND sg13g2_decap_8
XFILLER_122_147 VPWR VGND sg13g2_decap_8
XFILLER_104_840 VPWR VGND sg13g2_decap_8
X_12091_ VPWR _05937_ _05936_ VGND sg13g2_inv_1
XFILLER_1_422 VPWR VGND sg13g2_decap_8
XFILLER_110_309 VPWR VGND sg13g2_decap_8
X_11042_ acc_sum.exp_mant_logic0.a\[7\] _03343_ _05021_ VPWR VGND sg13g2_nor2_2
XFILLER_2_989 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_1_499 VPWR VGND sg13g2_decap_8
X_14801_ _00602_ VGND VPWR _01325_ acc_sum.exp_mant_logic0.a\[14\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
X_12993_ VPWR _06761_ _06760_ VGND sg13g2_inv_1
XFILLER_45_621 VPWR VGND sg13g2_fill_2
XFILLER_18_835 VPWR VGND sg13g2_decap_8
XFILLER_73_952 VPWR VGND sg13g2_decap_8
X_11944_ _05806_ VPWR _00986_ VGND net1874 _05805_ sg13g2_o21ai_1
X_14732_ _00533_ VGND VPWR _01260_ fp16_res_pipe.add_renorm0.exp\[3\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_2
XFILLER_72_451 VPWR VGND sg13g2_decap_8
X_14663_ _00464_ VGND VPWR _01191_ fp16_res_pipe.op_sign_logic0.mantisa_b\[0\] clknet_leaf_142_clk
+ sg13g2_dfrbpq_1
XFILLER_17_367 VPWR VGND sg13g2_decap_4
X_11875_ fp16_sum_pipe.reg3en.q\[0\] _05524_ _05540_ _05765_ VPWR VGND sg13g2_nand3_1
X_13614_ VPWR _00165_ net118 VGND sg13g2_inv_1
X_10826_ _04838_ _04722_ _04734_ VPWR VGND sg13g2_nand2_1
XFILLER_32_326 VPWR VGND sg13g2_decap_4
X_14594_ _00395_ VGND VPWR _01126_ fp16_res_pipe.y\[5\] clknet_leaf_129_clk sg13g2_dfrbpq_2
X_13545_ VPWR _00096_ net88 VGND sg13g2_inv_1
X_10757_ _04770_ _04733_ _04769_ VPWR VGND sg13g2_nand2_1
X_13476_ VPWR _00027_ net32 VGND sg13g2_inv_1
X_10688_ _04701_ _04700_ net1822 VPWR VGND sg13g2_nand2_1
XFILLER_127_932 VPWR VGND sg13g2_decap_8
X_12427_ VPWR VGND _06271_ _06272_ _06269_ _05997_ _06273_ _06268_ sg13g2_a221oi_1
XFILLER_9_599 VPWR VGND sg13g2_decap_8
XFILLER_126_475 VPWR VGND sg13g2_fill_2
XFILLER_114_626 VPWR VGND sg13g2_decap_8
X_12358_ _06190_ _06194_ _06203_ _06204_ VPWR VGND sg13g2_a21o_1
XFILLER_113_147 VPWR VGND sg13g2_fill_1
X_12289_ _06114_ _06134_ _06135_ VPWR VGND sg13g2_nor2_1
X_11309_ _05266_ net1812 _05161_ _05253_ net1654 VPWR VGND sg13g2_a22oi_1
XFILLER_45_1011 VPWR VGND sg13g2_fill_2
X_14028_ VPWR _00579_ net98 VGND sg13g2_inv_1
XFILLER_68_702 VPWR VGND sg13g2_decap_8
XFILLER_110_843 VPWR VGND sg13g2_decap_8
XFILLER_67_234 VPWR VGND sg13g2_decap_8
XFILLER_49_971 VPWR VGND sg13g2_fill_2
XFILLER_55_429 VPWR VGND sg13g2_fill_1
XFILLER_55_418 VPWR VGND sg13g2_decap_8
XFILLER_36_621 VPWR VGND sg13g2_fill_2
XFILLER_36_610 VPWR VGND sg13g2_fill_2
X_08520_ VPWR _02744_ _02743_ VGND sg13g2_inv_1
XFILLER_48_492 VPWR VGND sg13g2_decap_8
X_08451_ _02685_ _02683_ _02684_ VPWR VGND sg13g2_nand2_1
XFILLER_91_771 VPWR VGND sg13g2_decap_8
XFILLER_36_676 VPWR VGND sg13g2_decap_8
XFILLER_35_142 VPWR VGND sg13g2_fill_1
XFILLER_24_838 VPWR VGND sg13g2_decap_8
X_07402_ _01743_ acc_sub.exp_mant_logic0.a\[5\] VPWR VGND sg13g2_inv_2
XFILLER_63_495 VPWR VGND sg13g2_decap_8
XFILLER_51_657 VPWR VGND sg13g2_decap_8
XFILLER_51_635 VPWR VGND sg13g2_fill_2
XFILLER_50_112 VPWR VGND sg13g2_decap_8
XFILLER_35_175 VPWR VGND sg13g2_decap_8
XFILLER_23_337 VPWR VGND sg13g2_decap_8
X_08382_ _02568_ _02619_ _07114_ VPWR VGND sg13g2_nor2_1
X_07333_ _01694_ _01564_ _01695_ VPWR VGND sg13g2_and2_1
Xclkbuf_leaf_124_clk clknet_5_12__leaf_clk clknet_leaf_124_clk VPWR VGND sg13g2_buf_8
X_07264_ _01590_ VPWR _01634_ VGND _01500_ _01633_ sg13g2_o21ai_1
XFILLER_109_409 VPWR VGND sg13g2_fill_2
XFILLER_118_943 VPWR VGND sg13g2_decap_8
X_09003_ _03189_ _03180_ _03188_ VPWR VGND sg13g2_nand2_1
X_07195_ VPWR _01567_ _01566_ VGND sg13g2_inv_1
XFILLER_117_453 VPWR VGND sg13g2_decap_8
XFILLER_105_626 VPWR VGND sg13g2_fill_1
XFILLER_104_103 VPWR VGND sg13g2_fill_2
XFILLER_120_618 VPWR VGND sg13g2_fill_2
XFILLER_120_607 VPWR VGND sg13g2_decap_8
X_09905_ _03999_ _04001_ _04002_ VPWR VGND sg13g2_nor2_1
XFILLER_116_68 VPWR VGND sg13g2_decap_8
XFILLER_113_681 VPWR VGND sg13g2_fill_2
XFILLER_101_832 VPWR VGND sg13g2_decap_4
XFILLER_76_39 VPWR VGND sg13g2_fill_1
X_09836_ net1664 _03853_ _03946_ _03947_ VPWR VGND sg13g2_nand3_1
XFILLER_100_353 VPWR VGND sg13g2_fill_2
XFILLER_86_576 VPWR VGND sg13g2_fill_2
XFILLER_46_407 VPWR VGND sg13g2_decap_8
X_09767_ _03883_ _03882_ _03867_ VPWR VGND sg13g2_nand2_1
XFILLER_73_226 VPWR VGND sg13g2_fill_1
XFILLER_46_429 VPWR VGND sg13g2_decap_4
X_08718_ acc_sum.add_renorm0.exp\[4\] acc_sum.seg_reg0.q\[26\] net1819 _01331_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_73_248 VPWR VGND sg13g2_fill_1
XFILLER_39_481 VPWR VGND sg13g2_decap_8
XFILLER_27_643 VPWR VGND sg13g2_fill_2
X_08649_ net1816 acc_sum.add_renorm0.mantisa\[9\] _02870_ VPWR VGND sg13g2_nor2_1
XFILLER_82_760 VPWR VGND sg13g2_fill_1
XFILLER_54_451 VPWR VGND sg13g2_decap_8
XFILLER_42_613 VPWR VGND sg13g2_decap_8
Xclkbuf_5_2__f_clk clknet_4_1_0_clk clknet_5_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_25_21 VPWR VGND sg13g2_decap_8
XFILLER_109_1005 VPWR VGND sg13g2_decap_8
XFILLER_42_646 VPWR VGND sg13g2_decap_8
XFILLER_41_112 VPWR VGND sg13g2_decap_8
XFILLER_26_197 VPWR VGND sg13g2_decap_8
X_11660_ _05565_ _05470_ _05465_ _05477_ _05442_ VPWR VGND sg13g2_a22oi_1
XFILLER_23_860 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_115_clk clknet_5_8__leaf_clk clknet_leaf_115_clk VPWR VGND sg13g2_buf_8
X_10611_ VPWR _04624_ _04623_ VGND sg13g2_inv_1
X_11591_ _05495_ _05496_ VPWR VGND sg13g2_inv_4
X_13330_ _07036_ net1724 fp16_res_pipe.x2\[12\] VPWR VGND sg13g2_nand2_1
X_10542_ _04580_ _04501_ net1849 VPWR VGND sg13g2_nand2_1
XFILLER_127_217 VPWR VGND sg13g2_decap_8
XFILLER_109_921 VPWR VGND sg13g2_decap_8
X_13261_ acc\[12\] _06982_ net1679 _00846_ VPWR VGND sg13g2_mux2_1
XFILLER_41_42 VPWR VGND sg13g2_decap_8
X_12212_ _06058_ _06053_ _06055_ VPWR VGND sg13g2_nand2b_1
X_10473_ net1847 fp16_sum_pipe.add_renorm0.mantisa\[10\] _04521_ VPWR VGND sg13g2_nor2_1
XFILLER_124_935 VPWR VGND sg13g2_decap_8
XFILLER_109_998 VPWR VGND sg13g2_decap_8
XFILLER_108_486 VPWR VGND sg13g2_decap_4
X_13192_ VPWR _06929_ sipo.shift_reg\[7\] VGND sg13g2_inv_1
XFILLER_123_445 VPWR VGND sg13g2_decap_8
XFILLER_123_434 VPWR VGND sg13g2_decap_8
X_12143_ VGND VPWR _05914_ _05917_ _05989_ _05988_ sg13g2_a21oi_1
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_2_731 VPWR VGND sg13g2_decap_4
X_12074_ _05920_ _05919_ _05916_ VPWR VGND sg13g2_nand2_1
XFILLER_110_139 VPWR VGND sg13g2_fill_2
XFILLER_96_329 VPWR VGND sg13g2_fill_2
XFILLER_77_532 VPWR VGND sg13g2_fill_2
X_11025_ acc_sum.exp_mant_logic0.a\[11\] _03335_ _05004_ VPWR VGND sg13g2_nor2_1
XFILLER_2_786 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_92_513 VPWR VGND sg13g2_decap_4
XFILLER_18_610 VPWR VGND sg13g2_fill_1
XFILLER_92_546 VPWR VGND sg13g2_fill_1
XFILLER_92_535 VPWR VGND sg13g2_fill_1
XFILLER_46_963 VPWR VGND sg13g2_fill_2
XFILLER_46_930 VPWR VGND sg13g2_decap_8
X_12976_ _06746_ _06745_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_18_665 VPWR VGND sg13g2_decap_8
X_14715_ _00516_ VGND VPWR _01243_ fp16_res_pipe.exp_mant_logic0.a\[2\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_72_270 VPWR VGND sg13g2_decap_4
X_11927_ VPWR _05795_ fpmul.seg_reg0.q\[37\] VGND sg13g2_inv_1
XFILLER_17_197 VPWR VGND sg13g2_decap_4
XFILLER_32_123 VPWR VGND sg13g2_decap_4
XFILLER_33_635 VPWR VGND sg13g2_decap_8
XFILLER_60_465 VPWR VGND sg13g2_decap_8
X_14646_ _00447_ VGND VPWR net1916 fp16_res_pipe.reg1en.q\[0\] clknet_leaf_2_clk sg13g2_dfrbpq_2
XFILLER_33_668 VPWR VGND sg13g2_decap_8
XFILLER_14_860 VPWR VGND sg13g2_decap_8
X_11858_ _05755_ _05536_ _05665_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_106_clk clknet_5_14__leaf_clk clknet_leaf_106_clk VPWR VGND sg13g2_buf_8
X_11789_ _05691_ VPWR _01026_ VGND _05680_ _05690_ sg13g2_o21ai_1
X_14577_ _00378_ VGND VPWR _01109_ fp16_sum_pipe.exp_mant_logic0.b\[4\] clknet_leaf_117_clk
+ sg13g2_dfrbpq_2
X_10809_ _04774_ _04820_ _04821_ VPWR VGND sg13g2_nor2_1
X_13528_ VPWR _00079_ net26 VGND sg13g2_inv_1
XFILLER_118_217 VPWR VGND sg13g2_decap_8
X_13459_ _07109_ net1752 sipo.shift_reg\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_115_935 VPWR VGND sg13g2_decap_8
XFILLER_126_294 VPWR VGND sg13g2_decap_8
XFILLER_5_591 VPWR VGND sg13g2_fill_2
XFILLER_114_478 VPWR VGND sg13g2_decap_8
X_07951_ _01391_ _02183_ _02225_ _02182_ net1775 VPWR VGND sg13g2_a22oi_1
XFILLER_114_489 VPWR VGND sg13g2_fill_2
XFILLER_87_329 VPWR VGND sg13g2_decap_8
XFILLER_68_521 VPWR VGND sg13g2_decap_8
XFILLER_96_852 VPWR VGND sg13g2_decap_8
X_07882_ _02168_ net1887 acc_sub.x2\[8\] VPWR VGND sg13g2_nand2_1
X_09621_ _03738_ _03710_ _03723_ VPWR VGND sg13g2_nand2b_1
XFILLER_95_362 VPWR VGND sg13g2_decap_8
XFILLER_28_407 VPWR VGND sg13g2_decap_4
X_09552_ VPWR _03669_ acc_sum.add_renorm0.mantisa\[1\] VGND sg13g2_inv_1
XFILLER_37_952 VPWR VGND sg13g2_decap_8
X_08503_ acc_sum.seg_reg1.q\[21\] net1816 _02728_ VPWR VGND sg13g2_nor2_1
XFILLER_102_59 VPWR VGND sg13g2_decap_8
XFILLER_64_793 VPWR VGND sg13g2_decap_8
XFILLER_52_933 VPWR VGND sg13g2_decap_8
XFILLER_36_473 VPWR VGND sg13g2_decap_8
XFILLER_24_646 VPWR VGND sg13g2_fill_1
X_09483_ _03606_ VPWR _01247_ VGND net1917 _03605_ sg13g2_o21ai_1
X_08434_ fpdiv.divider0.remainder_reg\[6\] _01770_ _02667_ _02668_ VPWR VGND sg13g2_a21o_1
XFILLER_52_977 VPWR VGND sg13g2_decap_4
XFILLER_51_454 VPWR VGND sg13g2_fill_2
XFILLER_51_443 VPWR VGND sg13g2_fill_1
XFILLER_24_657 VPWR VGND sg13g2_decap_8
X_08365_ VPWR _02608_ _02607_ VGND sg13g2_inv_1
XFILLER_23_167 VPWR VGND sg13g2_fill_2
XFILLER_23_178 VPWR VGND sg13g2_fill_1
X_07316_ _01679_ VPWR _01680_ VGND _01541_ _01678_ sg13g2_o21ai_1
XFILLER_109_206 VPWR VGND sg13g2_decap_4
X_08296_ _02460_ _02345_ _02543_ VPWR VGND sg13g2_nor2_1
XFILLER_20_863 VPWR VGND sg13g2_decap_4
XFILLER_20_885 VPWR VGND sg13g2_decap_8
XFILLER_118_740 VPWR VGND sg13g2_decap_8
X_07247_ _01618_ _01617_ _01496_ VPWR VGND sg13g2_nand2_1
Xclkbuf_4_2_0_clk clknet_0_clk clknet_4_2_0_clk VPWR VGND sg13g2_buf_8
X_07178_ VPWR _01550_ acc_sub.op_sign_logic0.mantisa_b\[1\] VGND sg13g2_inv_1
XFILLER_11_56 VPWR VGND sg13g2_decap_8
XFILLER_127_56 VPWR VGND sg13g2_decap_8
XFILLER_106_957 VPWR VGND sg13g2_decap_8
XFILLER_79_808 VPWR VGND sg13g2_decap_8
XFILLER_3_539 VPWR VGND sg13g2_decap_8
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_121_938 VPWR VGND sg13g2_decap_8
XFILLER_87_830 VPWR VGND sg13g2_decap_8
XFILLER_78_329 VPWR VGND sg13g2_fill_1
XFILLER_59_521 VPWR VGND sg13g2_decap_4
XFILLER_59_510 VPWR VGND sg13g2_fill_2
XFILLER_87_841 VPWR VGND sg13g2_fill_2
XFILLER_59_565 VPWR VGND sg13g2_decap_8
X_09819_ _03783_ _03931_ _03928_ _03932_ VPWR VGND sg13g2_nand3_1
XFILLER_46_204 VPWR VGND sg13g2_decap_8
XFILLER_19_429 VPWR VGND sg13g2_fill_1
XFILLER_74_546 VPWR VGND sg13g2_decap_8
X_12830_ _06611_ VPWR _06612_ VGND net1958 _06609_ sg13g2_o21ai_1
XFILLER_28_952 VPWR VGND sg13g2_decap_8
XFILLER_74_579 VPWR VGND sg13g2_decap_8
XFILLER_36_42 VPWR VGND sg13g2_decap_8
XFILLER_27_440 VPWR VGND sg13g2_fill_1
X_12761_ VPWR _06546_ net1941 VGND sg13g2_inv_1
XFILLER_55_782 VPWR VGND sg13g2_decap_8
XFILLER_27_473 VPWR VGND sg13g2_decap_8
X_14500_ _00301_ VGND VPWR _01036_ fpdiv.reg_b_out\[7\] clknet_leaf_54_clk sg13g2_dfrbpq_2
X_12692_ _06501_ VPWR _00934_ VGND _06499_ net1741 sg13g2_o21ai_1
XFILLER_14_134 VPWR VGND sg13g2_decap_4
X_11712_ _05616_ fp16_sum_pipe.add_renorm0.exp\[1\] _05615_ VPWR VGND sg13g2_xnor2_1
X_14431_ _00232_ VGND VPWR _00970_ fpmul.seg_reg0.q\[16\] clknet_leaf_95_clk sg13g2_dfrbpq_1
XFILLER_42_487 VPWR VGND sg13g2_fill_1
X_11643_ _05548_ _05530_ _05504_ VPWR VGND sg13g2_xnor2_1
X_14362_ _00163_ VGND VPWR _00904_ _00015_ clknet_leaf_87_clk sg13g2_dfrbpq_1
XFILLER_52_96 VPWR VGND sg13g2_fill_1
XFILLER_6_300 VPWR VGND sg13g2_decap_8
X_11574_ _05472_ _05478_ _05467_ _05479_ VPWR VGND sg13g2_nand3_1
X_14293_ _00094_ VGND VPWR _00837_ acc\[3\] clknet_leaf_47_clk sg13g2_dfrbpq_2
X_13313_ _07023_ net1729 acc_sum.y\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_7_867 VPWR VGND sg13g2_decap_8
X_10525_ _04566_ _04564_ _04565_ _04562_ net1737 VPWR VGND sg13g2_a22oi_1
XFILLER_11_896 VPWR VGND sg13g2_decap_8
XFILLER_124_710 VPWR VGND sg13g2_fill_2
XFILLER_109_762 VPWR VGND sg13g2_fill_1
X_13244_ _06969_ net1676 _06968_ VPWR VGND sg13g2_nand2_1
X_10456_ _04503_ _04410_ _04502_ _04504_ VPWR VGND _04444_ sg13g2_nand4_1
XFILLER_124_732 VPWR VGND sg13g2_decap_8
X_13175_ _06917_ VPWR _00867_ VGND _06916_ net1712 sg13g2_o21ai_1
XFILLER_123_231 VPWR VGND sg13g2_decap_8
X_12126_ _05964_ _05947_ _05972_ VPWR VGND sg13g2_nor2_1
X_10387_ VPWR _04437_ _04436_ VGND sg13g2_inv_1
XFILLER_35_7 VPWR VGND sg13g2_decap_8
XFILLER_120_960 VPWR VGND sg13g2_decap_8
XFILLER_77_60 VPWR VGND sg13g2_decap_8
X_12057_ _05903_ _05901_ _05902_ VPWR VGND sg13g2_nand2_1
XFILLER_93_833 VPWR VGND sg13g2_decap_8
XFILLER_93_800 VPWR VGND sg13g2_decap_8
X_11008_ _04990_ fp16_res_pipe.x2\[0\] net1929 VPWR VGND sg13g2_nand2_1
XFILLER_92_310 VPWR VGND sg13g2_fill_1
XFILLER_93_877 VPWR VGND sg13g2_decap_8
XFILLER_53_708 VPWR VGND sg13g2_decap_8
XFILLER_19_985 VPWR VGND sg13g2_decap_8
X_12959_ _06729_ _06728_ fp16_sum_pipe.reg1en.d\[0\] _06730_ VPWR VGND sg13g2_a21o_2
XFILLER_52_229 VPWR VGND sg13g2_decap_4
XFILLER_34_933 VPWR VGND sg13g2_decap_8
XFILLER_18_484 VPWR VGND sg13g2_fill_2
XFILLER_60_273 VPWR VGND sg13g2_decap_8
X_14629_ _00430_ VGND VPWR _01161_ fp16_sum_pipe.add_renorm0.mantisa\[0\] clknet_leaf_109_clk
+ sg13g2_dfrbpq_1
XFILLER_33_487 VPWR VGND sg13g2_fill_1
XFILLER_119_504 VPWR VGND sg13g2_decap_8
XFILLER_14_690 VPWR VGND sg13g2_decap_4
X_08150_ _02410_ _02408_ _02273_ VPWR VGND sg13g2_nand2_1
XFILLER_119_537 VPWR VGND sg13g2_decap_8
XFILLER_9_182 VPWR VGND sg13g2_decap_4
X_08081_ _02305_ _02346_ _02347_ VPWR VGND sg13g2_nor2b_2
XFILLER_61_0 VPWR VGND sg13g2_decap_8
XFILLER_115_732 VPWR VGND sg13g2_decap_8
XFILLER_114_242 VPWR VGND sg13g2_decap_8
X_08983_ _01719_ VPWR _03169_ VGND _01721_ _03168_ sg13g2_o21ai_1
X_07934_ fp16_sum_pipe.exp_mant_logic0.b\[9\] _02208_ _02209_ VPWR VGND sg13g2_nor2_1
XFILLER_111_971 VPWR VGND sg13g2_decap_8
X_07865_ _02159_ _02153_ _02158_ VPWR VGND sg13g2_nand2_1
XFILLER_69_885 VPWR VGND sg13g2_decap_8
XFILLER_29_705 VPWR VGND sg13g2_decap_8
XFILLER_113_14 VPWR VGND sg13g2_decap_8
XFILLER_110_470 VPWR VGND sg13g2_fill_1
X_09604_ net1804 _03718_ _03720_ _03721_ VPWR VGND sg13g2_nor3_1
XFILLER_95_192 VPWR VGND sg13g2_decap_8
XFILLER_29_749 VPWR VGND sg13g2_decap_4
X_07796_ _02073_ _01939_ _01905_ _02095_ VPWR VGND sg13g2_nor3_1
X_09535_ _03652_ _03650_ _03651_ VPWR VGND sg13g2_xnor2_1
XFILLER_73_29 VPWR VGND sg13g2_decap_8
X_09466_ VPWR _03595_ fp16_res_pipe.exp_mant_logic0.a\[11\] VGND sg13g2_inv_1
XFILLER_40_903 VPWR VGND sg13g2_fill_1
XFILLER_24_443 VPWR VGND sg13g2_decap_8
XFILLER_25_966 VPWR VGND sg13g2_decap_8
X_08417_ _01756_ _02650_ _02652_ VPWR VGND sg13g2_nor2_2
XFILLER_52_774 VPWR VGND sg13g2_decap_8
XFILLER_51_273 VPWR VGND sg13g2_fill_1
XFILLER_40_958 VPWR VGND sg13g2_decap_4
X_09397_ _03420_ _03491_ net1675 _03543_ VPWR VGND sg13g2_mux2_1
X_08348_ _02591_ _02572_ _02561_ VPWR VGND sg13g2_nand2_1
XFILLER_7_119 VPWR VGND sg13g2_decap_8
X_08279_ _02528_ fp16_sum_pipe.exp_mant_logic0.b\[0\] _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[3\]
+ net1778 VPWR VGND sg13g2_a22oi_1
X_11290_ _03331_ _03333_ _03329_ _05250_ VPWR VGND _03335_ sg13g2_nand4_1
X_10310_ _04372_ VPWR _01186_ VGND net1914 _04005_ sg13g2_o21ai_1
XFILLER_4_804 VPWR VGND sg13g2_decap_8
XFILLER_106_721 VPWR VGND sg13g2_fill_2
XFILLER_98_59 VPWR VGND sg13g2_decap_8
X_10241_ _04128_ net1745 _04195_ _04313_ VPWR VGND sg13g2_nand3_1
XFILLER_106_765 VPWR VGND sg13g2_decap_4
XFILLER_79_627 VPWR VGND sg13g2_decap_8
XFILLER_78_115 VPWR VGND sg13g2_fill_1
XFILLER_78_104 VPWR VGND sg13g2_decap_8
X_10172_ _04252_ _04247_ _04251_ VPWR VGND sg13g2_nand2_1
XFILLER_120_245 VPWR VGND sg13g2_decap_8
XFILLER_87_682 VPWR VGND sg13g2_decap_8
XFILLER_75_800 VPWR VGND sg13g2_fill_2
XFILLER_59_362 VPWR VGND sg13g2_fill_2
XFILLER_59_351 VPWR VGND sg13g2_decap_8
X_13931_ VPWR _00482_ net6 VGND sg13g2_inv_1
XFILLER_102_993 VPWR VGND sg13g2_decap_8
XFILLER_75_833 VPWR VGND sg13g2_decap_4
XFILLER_90_825 VPWR VGND sg13g2_decap_8
XFILLER_47_96 VPWR VGND sg13g2_decap_8
X_13862_ VPWR _00413_ net51 VGND sg13g2_inv_1
XFILLER_19_248 VPWR VGND sg13g2_decap_8
X_13793_ VPWR _00344_ net74 VGND sg13g2_inv_1
X_12813_ _06596_ net1909 fp16_res_pipe.y\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_63_51 VPWR VGND sg13g2_decap_8
X_12744_ fpmul.reg_b_out\[13\] fp16_res_pipe.x2\[13\] net1952 _00923_ VPWR VGND sg13g2_mux2_1
XFILLER_16_966 VPWR VGND sg13g2_decap_8
XFILLER_31_914 VPWR VGND sg13g2_decap_8
X_12675_ VPWR _06488_ div_result\[11\] VGND sg13g2_inv_1
XFILLER_63_95 VPWR VGND sg13g2_decap_8
XFILLER_15_498 VPWR VGND sg13g2_fill_1
X_14414_ _00215_ VGND VPWR _00953_ fpmul.reg_a_out\[11\] clknet_leaf_125_clk sg13g2_dfrbpq_2
XFILLER_8_35 VPWR VGND sg13g2_decap_8
X_11626_ _05502_ _05530_ _05528_ _05531_ VPWR VGND sg13g2_nand3_1
XFILLER_30_468 VPWR VGND sg13g2_fill_1
X_14345_ _00146_ VGND VPWR _00887_ fpmul.reg_p_out\[9\] clknet_leaf_95_clk sg13g2_dfrbpq_1
XFILLER_11_671 VPWR VGND sg13g2_fill_1
XFILLER_11_682 VPWR VGND sg13g2_decap_8
X_11557_ _05462_ _05457_ _05461_ VPWR VGND sg13g2_nand2_2
XFILLER_7_664 VPWR VGND sg13g2_decap_8
X_10508_ VGND VPWR _04431_ _04436_ _04551_ _04433_ sg13g2_a21oi_1
X_11488_ _05397_ fp16_res_pipe.x2\[3\] net1945 VPWR VGND sg13g2_nand2_1
X_14276_ _00077_ VGND VPWR _00827_ fp16_res_pipe.x2\[9\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_98_925 VPWR VGND sg13g2_decap_8
X_13227_ net1742 _06952_ VPWR VGND sg13g2_inv_4
X_10439_ _04487_ VPWR _04488_ VGND _04442_ _04486_ sg13g2_o21ai_1
XFILLER_124_584 VPWR VGND sg13g2_decap_8
XFILLER_112_724 VPWR VGND sg13g2_fill_2
XFILLER_112_713 VPWR VGND sg13g2_decap_8
XFILLER_69_126 VPWR VGND sg13g2_fill_1
XFILLER_112_768 VPWR VGND sg13g2_decap_8
XFILLER_111_223 VPWR VGND sg13g2_fill_1
X_13089_ VGND VPWR fpmul.seg_reg0.q\[16\] fpmul.seg_reg0.q\[15\] _06851_ fpmul.seg_reg0.q\[17\]
+ sg13g2_a21oi_1
X_12109_ _05955_ _05952_ _05954_ VPWR VGND sg13g2_nand2_1
XFILLER_66_822 VPWR VGND sg13g2_decap_8
XFILLER_66_811 VPWR VGND sg13g2_decap_8
XFILLER_84_129 VPWR VGND sg13g2_decap_8
XFILLER_65_310 VPWR VGND sg13g2_decap_8
X_07650_ _01962_ _01869_ net1649 net1685 acc_sub.exp_mant_logic0.a\[4\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_81_814 VPWR VGND sg13g2_decap_8
X_07581_ _01894_ VPWR _01895_ VGND net1687 _01876_ sg13g2_o21ai_1
XFILLER_80_346 VPWR VGND sg13g2_fill_2
X_09320_ _03473_ _03472_ _03383_ VPWR VGND sg13g2_nand2_1
XFILLER_18_281 VPWR VGND sg13g2_decap_8
X_09251_ VPWR _03405_ fp16_res_pipe.op_sign_logic0.mantisa_a\[2\] VGND sg13g2_inv_1
X_08202_ VPWR _02458_ fp16_sum_pipe.exp_mant_logic0.b\[5\] VGND sg13g2_inv_1
XFILLER_22_947 VPWR VGND sg13g2_decap_8
XFILLER_119_301 VPWR VGND sg13g2_decap_8
X_09182_ _03344_ VPWR _01286_ VGND net1898 _03343_ sg13g2_o21ai_1
X_08133_ _02267_ _02380_ _02394_ VPWR VGND sg13g2_nor2_1
X_08064_ _02223_ VPWR _02330_ VGND _02329_ _02305_ sg13g2_o21ai_1
XFILLER_108_14 VPWR VGND sg13g2_decap_8
Xplace1820 acc_sum.reg3en.q\[0\] net1820 VPWR VGND sg13g2_buf_2
XFILLER_49_1009 VPWR VGND sg13g2_decap_4
Xplace1853 fpmul.seg_reg0.q\[15\] net1853 VPWR VGND sg13g2_buf_2
Xplace1831 fp16_res_pipe.reg1en.q\[0\] net1831 VPWR VGND sg13g2_buf_2
Xplace1842 fp16_sum_pipe.exp_mant_logic0.b\[5\] net1842 VPWR VGND sg13g2_buf_2
XFILLER_103_724 VPWR VGND sg13g2_fill_2
XFILLER_102_201 VPWR VGND sg13g2_decap_8
XFILLER_89_958 VPWR VGND sg13g2_decap_8
Xplace1886 net1885 net1886 VPWR VGND sg13g2_buf_1
Xplace1897 acc_sum.reg1en.d\[0\] net1897 VPWR VGND sg13g2_buf_1
Xplace1875 fpmul.reg1en.q\[0\] net1875 VPWR VGND sg13g2_buf_2
Xplace1864 fpmul.reg_b_out\[5\] net1864 VPWR VGND sg13g2_buf_2
XFILLER_0_306 VPWR VGND sg13g2_decap_8
XFILLER_1_829 VPWR VGND sg13g2_decap_8
XFILLER_103_768 VPWR VGND sg13g2_decap_8
XFILLER_124_35 VPWR VGND sg13g2_decap_8
X_08966_ acc_sub.add_renorm0.exp\[6\] net1699 _03152_ VPWR VGND sg13g2_nor2_1
X_08897_ _03000_ _02967_ _03083_ _03084_ VPWR VGND sg13g2_nor3_1
XFILLER_97_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_95_clk clknet_5_13__leaf_clk clknet_leaf_95_clk VPWR VGND sg13g2_buf_8
XFILLER_57_855 VPWR VGND sg13g2_decap_8
XFILLER_56_310 VPWR VGND sg13g2_decap_8
XFILLER_29_524 VPWR VGND sg13g2_decap_8
X_07917_ VPWR _02192_ fp16_sum_pipe.exp_mant_logic0.a\[11\] VGND sg13g2_inv_1
X_07848_ _02143_ _02006_ net1795 VPWR VGND sg13g2_nand2_1
XFILLER_56_354 VPWR VGND sg13g2_fill_2
XFILLER_56_343 VPWR VGND sg13g2_decap_8
XFILLER_16_229 VPWR VGND sg13g2_decap_8
X_07779_ _02080_ acc_sub.exp_mant_logic0.b\[4\] net1669 acc_sub.op_sign_logic0.mantisa_b\[7\]
+ net1781 VPWR VGND sg13g2_a22oi_1
X_09518_ _03635_ _03634_ _03624_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_77 VPWR VGND sg13g2_decap_4
XFILLER_25_774 VPWR VGND sg13g2_fill_1
X_10790_ VGND VPWR _04801_ _04802_ _04800_ net1709 sg13g2_a21oi_2
XFILLER_40_733 VPWR VGND sg13g2_decap_8
XFILLER_13_947 VPWR VGND sg13g2_decap_8
XFILLER_24_295 VPWR VGND sg13g2_fill_2
X_09449_ _03585_ net1832 fp16_res_pipe.seg_reg0.q\[24\] VPWR VGND sg13g2_nand2_1
XFILLER_33_21 VPWR VGND sg13g2_decap_8
X_12460_ _06302_ net1870 _06297_ _06303_ VPWR VGND sg13g2_nand3_1
XFILLER_32_1013 VPWR VGND sg13g2_fill_1
X_11411_ _05351_ VPWR _01064_ VGND _05350_ net1706 sg13g2_o21ai_1
X_12391_ VPWR VGND _06230_ _06236_ _06232_ _06235_ _06237_ _06226_ sg13g2_a221oi_1
XFILLER_8_439 VPWR VGND sg13g2_decap_4
XFILLER_21_980 VPWR VGND sg13g2_decap_8
XFILLER_126_827 VPWR VGND sg13g2_decap_8
X_14130_ VPWR _00681_ net119 VGND sg13g2_inv_1
X_11342_ _05296_ acc_sum.exp_mant_logic0.b\[1\] net1681 acc_sum.op_sign_logic0.mantisa_b\[4\]
+ net1762 VPWR VGND sg13g2_a22oi_1
XFILLER_125_315 VPWR VGND sg13g2_decap_8
XFILLER_109_0 VPWR VGND sg13g2_decap_8
X_14061_ VPWR _00612_ net94 VGND sg13g2_inv_1
X_11273_ _05235_ _05141_ acc_sum.exp_mant_logic0.a\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_3_133 VPWR VGND sg13g2_decap_8
XFILLER_79_402 VPWR VGND sg13g2_fill_1
XFILLER_4_678 VPWR VGND sg13g2_fill_2
X_10224_ _04297_ _04190_ net1745 fp16_res_pipe.exp_mant_logic0.b\[3\] net1644 VPWR
+ VGND sg13g2_a22oi_1
X_10155_ _04235_ VPWR _04236_ VGND _03613_ _04233_ sg13g2_o21ai_1
XFILLER_95_939 VPWR VGND sg13g2_decap_8
XFILLER_58_73 VPWR VGND sg13g2_fill_2
XFILLER_0_884 VPWR VGND sg13g2_decap_8
X_14963_ _00764_ VGND VPWR _01483_ acc_sub.add_renorm0.mantisa\[7\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_2
XFILLER_102_790 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_86_clk clknet_5_25__leaf_clk clknet_leaf_86_clk VPWR VGND sg13g2_buf_8
XFILLER_47_310 VPWR VGND sg13g2_fill_1
X_10086_ _03607_ _04156_ _04171_ VPWR VGND sg13g2_nor2_1
X_14894_ _00695_ VGND VPWR _01414_ acc_sub.op_sign_logic0.mantisa_b\[4\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_2
XFILLER_48_877 VPWR VGND sg13g2_decap_8
X_13914_ VPWR _00465_ net5 VGND sg13g2_inv_1
XFILLER_75_696 VPWR VGND sg13g2_decap_4
XFILLER_74_173 VPWR VGND sg13g2_decap_4
XFILLER_63_847 VPWR VGND sg13g2_fill_2
X_13845_ VPWR _00396_ net31 VGND sg13g2_inv_1
X_13776_ VPWR _00327_ net139 VGND sg13g2_inv_1
X_10988_ _04980_ fp16_res_pipe.x2\[10\] net1931 VPWR VGND sg13g2_nand2_1
X_12727_ _06513_ VPWR _06532_ VGND net1734 _06531_ sg13g2_o21ai_1
XFILLER_70_390 VPWR VGND sg13g2_decap_8
XFILLER_15_295 VPWR VGND sg13g2_decap_4
X_12658_ VGND VPWR _06413_ _06411_ _06474_ _06473_ sg13g2_a21oi_1
X_11609_ _05514_ _05513_ net1836 VPWR VGND sg13g2_nand2_1
XFILLER_30_298 VPWR VGND sg13g2_fill_1
XFILLER_117_816 VPWR VGND sg13g2_decap_8
X_12589_ _06405_ _06386_ _06383_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_10_clk clknet_5_4__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
XFILLER_8_951 VPWR VGND sg13g2_decap_8
X_14328_ _00129_ VGND VPWR _00871_ piso.tx_active clknet_leaf_57_clk sg13g2_dfrbpq_1
XFILLER_116_359 VPWR VGND sg13g2_decap_8
X_14259_ _00060_ VGND VPWR _00810_ acc_sub.x2\[8\] clknet_leaf_15_clk sg13g2_dfrbpq_2
XFILLER_125_893 VPWR VGND sg13g2_decap_8
X_08820_ _02971_ _03006_ _02991_ _02998_ _03007_ VPWR VGND sg13g2_nor4_1
XFILLER_112_521 VPWR VGND sg13g2_fill_2
XFILLER_97_232 VPWR VGND sg13g2_decap_8
XFILLER_86_917 VPWR VGND sg13g2_decap_8
XFILLER_57_107 VPWR VGND sg13g2_fill_2
XFILLER_24_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_77_clk clknet_5_27__leaf_clk clknet_leaf_77_clk VPWR VGND sg13g2_buf_8
XFILLER_85_449 VPWR VGND sg13g2_decap_8
XFILLER_85_438 VPWR VGND sg13g2_fill_1
X_08751_ VPWR _02947_ acc_sum.exp_mant_logic0.a\[8\] VGND sg13g2_inv_1
XFILLER_39_833 VPWR VGND sg13g2_decap_4
X_07702_ VGND VPWR _01869_ _02006_ _02010_ _02009_ sg13g2_a21oi_1
XFILLER_94_961 VPWR VGND sg13g2_decap_8
X_08682_ _02898_ _02896_ _02897_ _02895_ net1739 VPWR VGND sg13g2_a22oi_1
XFILLER_54_814 VPWR VGND sg13g2_fill_2
XFILLER_54_803 VPWR VGND sg13g2_decap_8
XFILLER_93_460 VPWR VGND sg13g2_fill_2
XFILLER_38_387 VPWR VGND sg13g2_fill_1
XFILLER_38_365 VPWR VGND sg13g2_decap_8
XFILLER_26_516 VPWR VGND sg13g2_decap_4
XFILLER_26_538 VPWR VGND sg13g2_fill_2
XFILLER_80_132 VPWR VGND sg13g2_decap_8
X_07564_ _01877_ VPWR _01878_ VGND _01787_ _01876_ sg13g2_o21ai_1
XFILLER_53_368 VPWR VGND sg13g2_decap_4
XFILLER_0_91 VPWR VGND sg13g2_decap_8
X_07495_ _01812_ _01817_ _01818_ VPWR VGND sg13g2_nor2_1
X_09303_ VGND VPWR _03453_ _03456_ _03457_ _03361_ sg13g2_a21oi_1
XFILLER_16_1008 VPWR VGND sg13g2_decap_4
X_09234_ _03385_ _03387_ _03388_ VPWR VGND sg13g2_nor2_2
X_09165_ _03333_ acc_sum.exp_mant_logic0.b\[12\] VPWR VGND sg13g2_inv_2
XFILLER_119_35 VPWR VGND sg13g2_decap_8
X_08116_ _02305_ _02377_ _02378_ VPWR VGND sg13g2_nor2b_2
X_09096_ _03276_ _03278_ _03274_ _03279_ VPWR VGND sg13g2_nand3_1
XFILLER_119_175 VPWR VGND sg13g2_decap_8
XFILLER_107_359 VPWR VGND sg13g2_decap_8
XFILLER_102_7 VPWR VGND sg13g2_decap_8
X_08047_ _02312_ VPWR _02313_ VGND _02229_ net1692 sg13g2_o21ai_1
Xplace1672 _01847_ net1672 VPWR VGND sg13g2_buf_2
Xplace1650 _01935_ net1650 VPWR VGND sg13g2_buf_1
Xplace1661 _05146_ net1661 VPWR VGND sg13g2_buf_1
XFILLER_103_521 VPWR VGND sg13g2_fill_2
Xplace1694 net1693 net1694 VPWR VGND sg13g2_buf_2
Xplace1683 _04052_ net1683 VPWR VGND sg13g2_buf_2
XFILLER_103_565 VPWR VGND sg13g2_decap_8
XFILLER_95_27 VPWR VGND sg13g2_fill_1
XFILLER_95_16 VPWR VGND sg13g2_decap_8
X_09998_ VPWR _04086_ _04085_ VGND sg13g2_inv_1
XFILLER_0_147 VPWR VGND sg13g2_decap_8
X_08949_ _03136_ _03135_ VPWR VGND sg13g2_inv_2
XFILLER_95_49 VPWR VGND sg13g2_decap_8
XFILLER_69_490 VPWR VGND sg13g2_decap_8
XFILLER_28_21 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_68_clk clknet_5_28__leaf_clk clknet_leaf_68_clk VPWR VGND sg13g2_buf_8
XFILLER_85_950 VPWR VGND sg13g2_decap_8
XFILLER_56_140 VPWR VGND sg13g2_fill_2
X_11960_ VPWR _05817_ fpmul.seg_reg0.q\[26\] VGND sg13g2_inv_1
XFILLER_72_622 VPWR VGND sg13g2_fill_1
XFILLER_72_600 VPWR VGND sg13g2_fill_2
X_10911_ _04920_ _04919_ _04741_ VPWR VGND sg13g2_nand2_1
X_11891_ VGND VPWR fpdiv.divider0.counter\[0\] _05767_ _01009_ _05776_ sg13g2_a21oi_1
XFILLER_44_357 VPWR VGND sg13g2_fill_2
XFILLER_44_324 VPWR VGND sg13g2_fill_2
XFILLER_71_165 VPWR VGND sg13g2_fill_2
XFILLER_60_828 VPWR VGND sg13g2_decap_8
X_13630_ VPWR _00181_ net29 VGND sg13g2_inv_1
XFILLER_44_42 VPWR VGND sg13g2_decap_8
X_10842_ _04784_ _04818_ _04851_ _04854_ VPWR VGND sg13g2_nand3_1
XFILLER_32_519 VPWR VGND sg13g2_decap_4
X_13561_ VPWR _00112_ net86 VGND sg13g2_inv_1
XFILLER_25_582 VPWR VGND sg13g2_decap_8
X_10773_ _04785_ _04784_ VPWR VGND sg13g2_inv_2
X_12512_ VPWR _06341_ acc_sub.x2\[10\] VGND sg13g2_inv_1
XFILLER_40_563 VPWR VGND sg13g2_decap_8
XFILLER_8_203 VPWR VGND sg13g2_decap_8
XFILLER_13_766 VPWR VGND sg13g2_fill_2
X_13492_ VPWR _00043_ net82 VGND sg13g2_inv_1
X_12443_ _06289_ _06283_ _06288_ VPWR VGND sg13g2_nand2_1
XFILLER_126_646 VPWR VGND sg13g2_decap_8
XFILLER_125_112 VPWR VGND sg13g2_decap_8
X_12374_ VGND VPWR _06220_ _06215_ _06214_ sg13g2_or2_1
X_11325_ _05277_ _05278_ _05279_ _05280_ VPWR VGND sg13g2_nor3_1
X_14113_ VPWR _00664_ net52 VGND sg13g2_inv_1
XFILLER_5_976 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_4_420 VPWR VGND sg13g2_decap_8
XFILLER_125_189 VPWR VGND sg13g2_decap_8
X_14044_ VPWR _00595_ net78 VGND sg13g2_inv_1
X_11256_ _01087_ _05218_ _05219_ VPWR VGND sg13g2_nand2_1
XFILLER_68_906 VPWR VGND sg13g2_fill_1
XFILLER_4_497 VPWR VGND sg13g2_decap_8
XFILLER_95_725 VPWR VGND sg13g2_fill_2
XFILLER_79_265 VPWR VGND sg13g2_decap_8
X_11187_ _05156_ _05075_ net1809 VPWR VGND sg13g2_nand2_1
XFILLER_69_94 VPWR VGND sg13g2_fill_1
X_10207_ _04282_ net1829 net1643 net1688 fp16_res_pipe.exp_mant_logic0.b\[4\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_122_896 VPWR VGND sg13g2_decap_8
XFILLER_121_395 VPWR VGND sg13g2_fill_1
XFILLER_121_384 VPWR VGND sg13g2_decap_4
XFILLER_48_630 VPWR VGND sg13g2_fill_1
X_10138_ _04220_ _04219_ _04150_ VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_59_clk clknet_5_30__leaf_clk clknet_leaf_59_clk VPWR VGND sg13g2_buf_8
XFILLER_95_769 VPWR VGND sg13g2_decap_4
X_14946_ _00747_ VGND VPWR _01466_ acc_sub.exp_mant_logic0.a\[14\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_1
XFILLER_85_60 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_fill_1
X_10069_ _04156_ net1662 _04144_ VPWR VGND sg13g2_nand2_2
XFILLER_78_1013 VPWR VGND sg13g2_fill_1
XFILLER_36_836 VPWR VGND sg13g2_fill_2
X_14877_ _00678_ VGND VPWR _01397_ acc_sub.exp_mant_logic0.b\[3\] clknet_leaf_59_clk
+ sg13g2_dfrbpq_2
XFILLER_62_132 VPWR VGND sg13g2_decap_8
XFILLER_35_324 VPWR VGND sg13g2_decap_8
XFILLER_91_975 VPWR VGND sg13g2_decap_8
XFILLER_62_165 VPWR VGND sg13g2_fill_1
XFILLER_50_305 VPWR VGND sg13g2_decap_8
X_13828_ VPWR _00379_ net47 VGND sg13g2_inv_1
X_13759_ VPWR _00310_ net129 VGND sg13g2_inv_1
X_07280_ _01508_ _01611_ _01648_ VPWR VGND sg13g2_nor2_1
XFILLER_31_530 VPWR VGND sg13g2_decap_4
XFILLER_31_541 VPWR VGND sg13g2_fill_1
XFILLER_31_552 VPWR VGND sg13g2_fill_1
XFILLER_102_1000 VPWR VGND sg13g2_decap_8
XFILLER_116_145 VPWR VGND sg13g2_decap_8
XFILLER_85_1006 VPWR VGND sg13g2_decap_8
XFILLER_7_291 VPWR VGND sg13g2_decap_8
XFILLER_104_329 VPWR VGND sg13g2_decap_8
X_09921_ VPWR _04018_ fp16_res_pipe.exp_mant_logic0.b\[10\] VGND sg13g2_inv_1
XFILLER_113_830 VPWR VGND sg13g2_decap_8
XFILLER_98_541 VPWR VGND sg13g2_decap_4
XFILLER_98_530 VPWR VGND sg13g2_fill_2
XFILLER_112_351 VPWR VGND sg13g2_decap_8
X_09852_ _03962_ _03846_ _03845_ VPWR VGND sg13g2_nand2_1
XFILLER_105_15 VPWR VGND sg13g2_decap_8
XFILLER_98_563 VPWR VGND sg13g2_decap_8
X_08803_ _02990_ _02981_ _02989_ VPWR VGND sg13g2_nand2_2
X_09783_ VPWR _03898_ _03823_ VGND sg13g2_inv_1
XFILLER_98_596 VPWR VGND sg13g2_fill_1
XFILLER_98_585 VPWR VGND sg13g2_decap_8
XFILLER_85_257 VPWR VGND sg13g2_decap_8
X_08734_ _02936_ acc\[14\] net1901 VPWR VGND sg13g2_nand2_1
XFILLER_27_803 VPWR VGND sg13g2_fill_2
XFILLER_94_780 VPWR VGND sg13g2_fill_1
XFILLER_38_140 VPWR VGND sg13g2_fill_2
XFILLER_27_825 VPWR VGND sg13g2_decap_8
XFILLER_121_14 VPWR VGND sg13g2_decap_8
X_08665_ VGND VPWR _02882_ net1818 _01342_ _02883_ sg13g2_a21oi_1
XFILLER_93_290 VPWR VGND sg13g2_decap_4
XFILLER_82_975 VPWR VGND sg13g2_decap_8
X_08596_ _02819_ acc_sum.op_sign_logic0.mantisa_a\[1\] acc_sum.op_sign_logic0.mantisa_b\[1\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_42_817 VPWR VGND sg13g2_decap_8
X_07547_ _01863_ acc_sub.exp_mant_logic0.a\[7\] _01847_ _01779_ acc_sub.seg_reg0.q\[22\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_81_485 VPWR VGND sg13g2_decap_8
XFILLER_22_541 VPWR VGND sg13g2_fill_1
X_07478_ _01798_ _01800_ _01801_ VPWR VGND sg13g2_nor2_1
XFILLER_50_894 VPWR VGND sg13g2_decap_8
XFILLER_14_56 VPWR VGND sg13g2_decap_8
XFILLER_6_707 VPWR VGND sg13g2_decap_8
X_09217_ fp16_res_pipe.op_sign_logic0.mantisa_b\[8\] _03370_ _03371_ VPWR VGND sg13g2_nor2_1
XFILLER_14_89 VPWR VGND sg13g2_fill_2
XFILLER_108_613 VPWR VGND sg13g2_decap_8
XFILLER_107_112 VPWR VGND sg13g2_decap_8
X_09148_ acc_sub.reg3en.q\[0\] acc_sub.y\[3\] _03323_ VPWR VGND sg13g2_nor2_1
XFILLER_5_206 VPWR VGND sg13g2_fill_1
X_09079_ _03262_ _03183_ _03263_ VPWR VGND sg13g2_nor2b_1
XFILLER_108_668 VPWR VGND sg13g2_decap_8
XFILLER_107_156 VPWR VGND sg13g2_decap_4
XFILLER_100_4 VPWR VGND sg13g2_fill_1
X_11110_ _05018_ _05079_ _05080_ VPWR VGND sg13g2_nor2_1
XFILLER_1_401 VPWR VGND sg13g2_decap_8
XFILLER_30_77 VPWR VGND sg13g2_decap_8
XFILLER_122_126 VPWR VGND sg13g2_decap_8
X_12090_ _05936_ net1867 _05935_ VPWR VGND sg13g2_xnor2_1
X_11041_ VPWR _05020_ _05019_ VGND sg13g2_inv_1
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_2_968 VPWR VGND sg13g2_decap_8
XFILLER_103_362 VPWR VGND sg13g2_fill_2
XFILLER_89_585 VPWR VGND sg13g2_decap_4
XFILLER_77_758 VPWR VGND sg13g2_fill_2
XFILLER_77_725 VPWR VGND sg13g2_decap_8
XFILLER_76_213 VPWR VGND sg13g2_fill_1
XFILLER_49_416 VPWR VGND sg13g2_decap_8
XFILLER_1_478 VPWR VGND sg13g2_decap_8
XFILLER_76_268 VPWR VGND sg13g2_fill_2
XFILLER_65_909 VPWR VGND sg13g2_fill_1
X_14800_ _00601_ VGND VPWR _01324_ acc_sum.exp_mant_logic0.a\[13\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
XFILLER_58_950 VPWR VGND sg13g2_decap_8
X_12992_ _06760_ fpmul.seg_reg0.q\[19\] _06752_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_313 VPWR VGND sg13g2_fill_1
XFILLER_29_162 VPWR VGND sg13g2_fill_2
XFILLER_72_430 VPWR VGND sg13g2_decap_8
XFILLER_57_493 VPWR VGND sg13g2_fill_2
X_11943_ _05806_ net1874 fpmul.reg_b_out\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_18_858 VPWR VGND sg13g2_fill_2
X_14731_ _00532_ VGND VPWR _01259_ fp16_res_pipe.add_renorm0.exp\[2\] clknet_leaf_132_clk
+ sg13g2_dfrbpq_1
XFILLER_44_154 VPWR VGND sg13g2_fill_2
X_11874_ VPWR _05764_ add_result\[0\] VGND sg13g2_inv_1
X_14662_ _00463_ VGND VPWR _01190_ fp16_res_pipe.exp_mant_logic0.b\[15\] clknet_leaf_130_clk
+ sg13g2_dfrbpq_1
XFILLER_33_806 VPWR VGND sg13g2_decap_8
X_13613_ VPWR _00164_ net112 VGND sg13g2_inv_1
XFILLER_60_647 VPWR VGND sg13g2_fill_1
X_10825_ _04837_ _04824_ VPWR VGND sg13g2_inv_2
XFILLER_26_891 VPWR VGND sg13g2_decap_8
XFILLER_111_91 VPWR VGND sg13g2_decap_8
X_14593_ _00394_ VGND VPWR _01125_ fp16_res_pipe.y\[4\] clknet_leaf_127_clk sg13g2_dfrbpq_1
XFILLER_32_349 VPWR VGND sg13g2_decap_8
X_13544_ VPWR _00095_ net100 VGND sg13g2_inv_1
XFILLER_41_872 VPWR VGND sg13g2_fill_1
X_10756_ _04745_ _04755_ _04760_ _04768_ _04769_ VPWR VGND sg13g2_nor4_1
XFILLER_127_911 VPWR VGND sg13g2_decap_8
X_13475_ VPWR _00026_ net33 VGND sg13g2_inv_1
XFILLER_40_382 VPWR VGND sg13g2_decap_8
X_10687_ _04697_ _04698_ _04696_ _04700_ VPWR VGND _04699_ sg13g2_nand4_1
XFILLER_65_7 VPWR VGND sg13g2_fill_2
X_12426_ _06257_ _06256_ _06272_ VPWR VGND sg13g2_nor2b_1
XFILLER_127_988 VPWR VGND sg13g2_decap_8
X_12357_ _06015_ _06165_ _06192_ _06203_ VPWR VGND sg13g2_nor3_1
XFILLER_5_773 VPWR VGND sg13g2_decap_8
XFILLER_113_126 VPWR VGND sg13g2_decap_8
X_12288_ _06134_ _06131_ _06133_ VPWR VGND sg13g2_nand2_1
X_11308_ _01081_ _05264_ _05265_ VPWR VGND sg13g2_nand2_1
X_14027_ VPWR _00578_ net103 VGND sg13g2_inv_1
XFILLER_95_500 VPWR VGND sg13g2_decap_8
X_11239_ _05203_ net1661 net1810 VPWR VGND sg13g2_nand2_1
XFILLER_110_822 VPWR VGND sg13g2_decap_8
XFILLER_96_70 VPWR VGND sg13g2_decap_8
XFILLER_1_990 VPWR VGND sg13g2_decap_8
XFILLER_110_899 VPWR VGND sg13g2_decap_8
XFILLER_64_920 VPWR VGND sg13g2_decap_8
X_14929_ _00730_ VGND VPWR _01449_ fpdiv.divider0.divisor_reg\[9\] clknet_leaf_75_clk
+ sg13g2_dfrbpq_2
XFILLER_82_249 VPWR VGND sg13g2_decap_8
XFILLER_36_633 VPWR VGND sg13g2_fill_1
X_08450_ VPWR _02684_ fpdiv.divider0.remainder_reg\[12\] VGND sg13g2_inv_1
XFILLER_64_975 VPWR VGND sg13g2_decap_8
XFILLER_63_441 VPWR VGND sg13g2_fill_1
XFILLER_24_806 VPWR VGND sg13g2_decap_8
XFILLER_24_817 VPWR VGND sg13g2_fill_2
XFILLER_91_1010 VPWR VGND sg13g2_decap_4
X_07401_ _01742_ VPWR _01458_ VGND net1890 _01741_ sg13g2_o21ai_1
X_08381_ _02621_ _07116_ fpmul.reg3en.q\[0\] VPWR VGND sg13g2_nand2b_1
XFILLER_17_891 VPWR VGND sg13g2_decap_8
XFILLER_23_316 VPWR VGND sg13g2_decap_8
X_07332_ _01693_ VPWR _01694_ VGND _01553_ net1666 sg13g2_o21ai_1
XFILLER_91_0 VPWR VGND sg13g2_decap_8
XFILLER_50_168 VPWR VGND sg13g2_decap_8
XFILLER_32_883 VPWR VGND sg13g2_fill_2
XFILLER_32_894 VPWR VGND sg13g2_decap_8
X_07263_ VPWR VGND _01515_ _01512_ _01632_ _01506_ _01633_ _01513_ sg13g2_a221oi_1
X_07194_ _01559_ _01565_ _01566_ VPWR VGND sg13g2_nor2_1
XFILLER_118_922 VPWR VGND sg13g2_decap_8
XFILLER_117_410 VPWR VGND sg13g2_decap_4
X_09002_ _03183_ _03187_ _03188_ VPWR VGND sg13g2_nor2_1
XFILLER_117_432 VPWR VGND sg13g2_decap_8
XFILLER_118_999 VPWR VGND sg13g2_decap_8
XFILLER_105_649 VPWR VGND sg13g2_decap_4
XFILLER_104_137 VPWR VGND sg13g2_decap_8
XFILLER_116_47 VPWR VGND sg13g2_decap_8
XFILLER_104_148 VPWR VGND sg13g2_fill_2
X_09904_ fp16_res_pipe.exp_mant_logic0.a\[13\] _04000_ _04001_ VPWR VGND sg13g2_nor2_1
XFILLER_113_693 VPWR VGND sg13g2_fill_1
X_09835_ _03843_ _03847_ _03852_ _03946_ VPWR VGND sg13g2_or3_1
XFILLER_101_811 VPWR VGND sg13g2_decap_8
XFILLER_101_866 VPWR VGND sg13g2_decap_8
XFILLER_100_321 VPWR VGND sg13g2_decap_8
XFILLER_86_555 VPWR VGND sg13g2_decap_8
X_09766_ _03838_ _03881_ _03882_ VPWR VGND sg13g2_nor2_2
XFILLER_101_899 VPWR VGND sg13g2_decap_8
XFILLER_86_588 VPWR VGND sg13g2_decap_8
XFILLER_74_739 VPWR VGND sg13g2_decap_8
X_09697_ _03809_ _03812_ _03813_ VPWR VGND sg13g2_and2_1
X_08717_ _02925_ VPWR _01332_ VGND net1814 _02924_ sg13g2_o21ai_1
XFILLER_55_942 VPWR VGND sg13g2_decap_8
XFILLER_27_633 VPWR VGND sg13g2_fill_2
X_08648_ _02869_ _02788_ _02868_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_666 VPWR VGND sg13g2_decap_4
XFILLER_26_187 VPWR VGND sg13g2_fill_1
X_08579_ _02803_ acc_sum.reg2en.q\[0\] VPWR VGND sg13g2_inv_2
XFILLER_70_978 VPWR VGND sg13g2_decap_4
XFILLER_23_850 VPWR VGND sg13g2_decap_4
X_10610_ _04622_ VPWR _04623_ VGND net1826 fp16_res_pipe.add_renorm0.mantisa\[4\]
+ sg13g2_o21ai_1
X_11590_ _05475_ _05494_ _05495_ VPWR VGND sg13g2_nor2_2
XFILLER_109_900 VPWR VGND sg13g2_decap_8
XFILLER_41_21 VPWR VGND sg13g2_decap_8
X_10541_ VPWR _04579_ fp16_sum_pipe.add_renorm0.mantisa\[0\] VGND sg13g2_inv_1
X_13260_ _06981_ VPWR _06982_ VGND _06980_ _06952_ sg13g2_o21ai_1
XFILLER_109_977 VPWR VGND sg13g2_decap_8
XFILLER_108_443 VPWR VGND sg13g2_fill_2
XFILLER_108_432 VPWR VGND sg13g2_decap_8
XFILLER_68_1012 VPWR VGND sg13g2_fill_2
X_12211_ VPWR _06057_ _06056_ VGND sg13g2_inv_1
XFILLER_41_98 VPWR VGND sg13g2_decap_8
XFILLER_6_537 VPWR VGND sg13g2_fill_2
X_10472_ _04520_ _04499_ _04519_ VPWR VGND sg13g2_xnor2_1
XFILLER_124_914 VPWR VGND sg13g2_decap_8
X_13191_ _06928_ VPWR _00862_ VGND _06927_ net1712 sg13g2_o21ai_1
XFILLER_97_809 VPWR VGND sg13g2_fill_2
X_12142_ VPWR _05988_ _05915_ VGND sg13g2_inv_1
XFILLER_123_479 VPWR VGND sg13g2_decap_8
X_12073_ _05919_ _05914_ _05915_ VPWR VGND sg13g2_nand2_1
XFILLER_89_371 VPWR VGND sg13g2_decap_8
XFILLER_77_511 VPWR VGND sg13g2_decap_8
X_11024_ acc_sum.exp_mant_logic0.b\[11\] _02941_ _05003_ VPWR VGND sg13g2_nor2_1
XFILLER_49_213 VPWR VGND sg13g2_decap_8
XFILLER_77_544 VPWR VGND sg13g2_decap_8
XFILLER_77_588 VPWR VGND sg13g2_decap_8
XFILLER_49_279 VPWR VGND sg13g2_decap_8
XFILLER_46_920 VPWR VGND sg13g2_decap_4
XFILLER_37_419 VPWR VGND sg13g2_fill_2
XFILLER_37_408 VPWR VGND sg13g2_decap_8
X_12975_ _06744_ VPWR _06745_ VGND net1962 _06742_ sg13g2_o21ai_1
XFILLER_66_95 VPWR VGND sg13g2_decap_4
XFILLER_57_290 VPWR VGND sg13g2_fill_2
XFILLER_73_772 VPWR VGND sg13g2_decap_8
XFILLER_73_761 VPWR VGND sg13g2_fill_2
XFILLER_73_750 VPWR VGND sg13g2_decap_8
X_11926_ _05794_ VPWR _00992_ VGND net1879 _05793_ sg13g2_o21ai_1
X_14714_ _00515_ VGND VPWR _01242_ fp16_res_pipe.exp_mant_logic0.a\[1\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
XFILLER_61_945 VPWR VGND sg13g2_decap_4
XFILLER_17_165 VPWR VGND sg13g2_decap_4
XFILLER_32_113 VPWR VGND sg13g2_fill_1
XFILLER_33_614 VPWR VGND sg13g2_decap_8
XFILLER_82_83 VPWR VGND sg13g2_decap_4
XFILLER_61_989 VPWR VGND sg13g2_fill_2
X_14645_ _00446_ VGND VPWR fp16_res_pipe.reg1en.q\[0\] fp16_res_pipe.reg2en.q\[0\]
+ clknet_leaf_139_clk sg13g2_dfrbpq_2
X_11857_ _05754_ _05537_ _05665_ VPWR VGND sg13g2_nand2b_1
X_11788_ _05691_ _05573_ add_result\[13\] VPWR VGND sg13g2_nand2_1
X_14576_ _00377_ VGND VPWR _01108_ fp16_sum_pipe.exp_mant_logic0.b\[3\] clknet_leaf_135_clk
+ sg13g2_dfrbpq_2
XFILLER_32_179 VPWR VGND sg13g2_decap_8
X_10808_ _04820_ _04785_ _04819_ VPWR VGND sg13g2_xnor2_1
X_13527_ VPWR _00078_ net35 VGND sg13g2_inv_1
X_10739_ _04750_ _04636_ _04752_ VPWR VGND sg13g2_and2_1
X_13458_ _07108_ VPWR _00775_ VGND _06931_ net1752 sg13g2_o21ai_1
XFILLER_127_785 VPWR VGND sg13g2_decap_8
XFILLER_115_914 VPWR VGND sg13g2_decap_8
XFILLER_114_402 VPWR VGND sg13g2_fill_2
X_13389_ acc_sub.x2\[4\] net1693 _07071_ VPWR VGND sg13g2_nor2_1
X_12409_ _06255_ _05781_ _06254_ VPWR VGND sg13g2_xnor2_1
XFILLER_126_273 VPWR VGND sg13g2_decap_8
XFILLER_114_424 VPWR VGND sg13g2_decap_8
XFILLER_99_146 VPWR VGND sg13g2_decap_8
X_07950_ _02225_ _02223_ fp16_sum_pipe.exp_mant_logic0.a\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_68_500 VPWR VGND sg13g2_decap_8
X_07881_ _02167_ VPWR _01403_ VGND net1895 _01808_ sg13g2_o21ai_1
XFILLER_95_330 VPWR VGND sg13g2_decap_4
XFILLER_56_706 VPWR VGND sg13g2_decap_8
X_09620_ _03737_ _03735_ _03714_ VPWR VGND sg13g2_nand2_1
XFILLER_55_205 VPWR VGND sg13g2_fill_1
XFILLER_83_558 VPWR VGND sg13g2_decap_4
XFILLER_55_249 VPWR VGND sg13g2_fill_2
XFILLER_49_780 VPWR VGND sg13g2_fill_2
XFILLER_37_931 VPWR VGND sg13g2_decap_8
XFILLER_64_772 VPWR VGND sg13g2_fill_2
XFILLER_64_761 VPWR VGND sg13g2_decap_4
XFILLER_64_783 VPWR VGND sg13g2_decap_4
XFILLER_51_422 VPWR VGND sg13g2_decap_4
XFILLER_24_636 VPWR VGND sg13g2_decap_4
X_09482_ _03606_ acc_sub.x2\[6\] net1916 VPWR VGND sg13g2_nand2_1
X_08433_ _02660_ _02666_ _02667_ VPWR VGND sg13g2_nor2_1
XFILLER_52_956 VPWR VGND sg13g2_decap_8
XFILLER_23_146 VPWR VGND sg13g2_fill_1
X_08364_ instr\[1\] instr\[0\] _02607_ VPWR VGND sg13g2_nor2_1
XFILLER_51_477 VPWR VGND sg13g2_fill_2
XFILLER_51_466 VPWR VGND sg13g2_decap_8
X_07315_ VGND VPWR _01678_ _01541_ _01679_ _01656_ sg13g2_a21oi_1
X_08295_ _02468_ _02349_ _02542_ VPWR VGND sg13g2_nor2_1
X_07246_ _01616_ VPWR _01617_ VGND _01499_ _01501_ sg13g2_o21ai_1
X_07177_ _01549_ _01548_ acc_sub.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_3_518 VPWR VGND sg13g2_decap_8
XFILLER_11_35 VPWR VGND sg13g2_decap_8
XFILLER_127_35 VPWR VGND sg13g2_decap_8
XFILLER_118_796 VPWR VGND sg13g2_decap_8
XFILLER_117_273 VPWR VGND sg13g2_decap_4
XFILLER_106_936 VPWR VGND sg13g2_decap_8
XFILLER_105_413 VPWR VGND sg13g2_decap_8
XFILLER_121_917 VPWR VGND sg13g2_decap_8
XFILLER_105_479 VPWR VGND sg13g2_decap_8
XFILLER_87_39 VPWR VGND sg13g2_decap_8
XFILLER_87_28 VPWR VGND sg13g2_fill_1
XFILLER_101_630 VPWR VGND sg13g2_fill_1
XFILLER_98_190 VPWR VGND sg13g2_decap_8
XFILLER_87_853 VPWR VGND sg13g2_fill_1
XFILLER_101_685 VPWR VGND sg13g2_decap_8
X_09818_ net1769 VPWR _03931_ VGND _03929_ _03930_ sg13g2_o21ai_1
XFILLER_100_140 VPWR VGND sg13g2_fill_1
XFILLER_87_886 VPWR VGND sg13g2_decap_8
XFILLER_86_374 VPWR VGND sg13g2_fill_2
X_09749_ _03865_ _03864_ VPWR VGND sg13g2_inv_2
XFILLER_36_21 VPWR VGND sg13g2_decap_8
XFILLER_28_931 VPWR VGND sg13g2_decap_8
XFILLER_62_709 VPWR VGND sg13g2_decap_4
XFILLER_43_901 VPWR VGND sg13g2_fill_1
XFILLER_61_219 VPWR VGND sg13g2_fill_1
X_12760_ fpmul.reg_b_out\[0\] fp16_res_pipe.x2\[0\] net1957 _00910_ VPWR VGND sg13g2_mux2_1
XFILLER_82_591 VPWR VGND sg13g2_fill_1
X_12691_ _06479_ VPWR _06501_ VGND net1734 _06500_ sg13g2_o21ai_1
XFILLER_36_98 VPWR VGND sg13g2_decap_8
XFILLER_14_124 VPWR VGND sg13g2_fill_2
X_11711_ _05615_ _05583_ fp16_sum_pipe.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
X_14430_ _00231_ VGND VPWR _00969_ fpmul.seg_reg0.q\[15\] clknet_leaf_101_clk sg13g2_dfrbpq_2
XFILLER_14_179 VPWR VGND sg13g2_fill_2
X_11642_ net1836 VPWR _05547_ VGND _05542_ _05546_ sg13g2_o21ai_1
XFILLER_30_628 VPWR VGND sg13g2_decap_4
X_14361_ _00162_ VGND VPWR _00903_ _00014_ clknet_leaf_87_clk sg13g2_dfrbpq_1
XFILLER_23_691 VPWR VGND sg13g2_decap_4
X_13312_ _07022_ _02578_ acc_sub.y\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_11_875 VPWR VGND sg13g2_decap_8
X_11573_ _05478_ _05475_ _05477_ VPWR VGND sg13g2_nand2_1
X_14292_ _00093_ VGND VPWR _00836_ acc\[2\] clknet_leaf_45_clk sg13g2_dfrbpq_2
XFILLER_7_846 VPWR VGND sg13g2_decap_8
X_10524_ VGND VPWR net1670 _04508_ _04565_ net1737 sg13g2_a21oi_1
X_13243_ _06966_ _06967_ _06965_ _06968_ VPWR VGND sg13g2_nand3_1
X_10455_ _04499_ _04451_ _04454_ _04503_ VPWR VGND sg13g2_nor3_1
XFILLER_123_210 VPWR VGND sg13g2_decap_8
X_13174_ _06917_ net1712 sipo.word\[12\] VPWR VGND sg13g2_nand2_1
X_12125_ _05970_ _05966_ _05971_ VPWR VGND sg13g2_xor2_1
X_10386_ _04433_ _04435_ _04436_ VPWR VGND sg13g2_nor2_2
XFILLER_2_551 VPWR VGND sg13g2_fill_1
XFILLER_124_788 VPWR VGND sg13g2_decap_8
XFILLER_123_287 VPWR VGND sg13g2_decap_8
X_12056_ _05902_ net1856 net1865 VPWR VGND sg13g2_nand2_1
XFILLER_42_1004 VPWR VGND sg13g2_decap_8
XFILLER_28_7 VPWR VGND sg13g2_decap_8
XFILLER_77_363 VPWR VGND sg13g2_fill_1
XFILLER_65_514 VPWR VGND sg13g2_decap_8
XFILLER_65_503 VPWR VGND sg13g2_decap_8
X_11007_ _04989_ VPWR _01106_ VGND net1928 _02460_ sg13g2_o21ai_1
XFILLER_92_322 VPWR VGND sg13g2_decap_8
XFILLER_92_366 VPWR VGND sg13g2_decap_8
XFILLER_80_506 VPWR VGND sg13g2_fill_2
XFILLER_65_569 VPWR VGND sg13g2_decap_8
XFILLER_18_452 VPWR VGND sg13g2_fill_1
XFILLER_19_964 VPWR VGND sg13g2_decap_8
X_12958_ _06729_ net1910 fp16_res_pipe.y\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_46_794 VPWR VGND sg13g2_decap_8
XFILLER_34_912 VPWR VGND sg13g2_decap_8
XFILLER_18_463 VPWR VGND sg13g2_decap_8
XFILLER_33_411 VPWR VGND sg13g2_fill_1
X_12889_ VPWR _06666_ fpmul.reg_p_out\[7\] VGND sg13g2_inv_1
X_11909_ _05783_ fpmul.reg_a_out\[4\] VPWR VGND sg13g2_inv_2
XFILLER_33_455 VPWR VGND sg13g2_decap_8
XFILLER_61_797 VPWR VGND sg13g2_decap_8
XFILLER_60_252 VPWR VGND sg13g2_decap_8
XFILLER_34_989 VPWR VGND sg13g2_decap_8
X_14628_ _00429_ VGND VPWR _01160_ fp16_sum_pipe.add_renorm0.exp\[7\] clknet_leaf_98_clk
+ sg13g2_dfrbpq_1
X_14559_ _00360_ VGND VPWR _01095_ acc_sum.seg_reg0.q\[22\] clknet_leaf_25_clk sg13g2_dfrbpq_1
XFILLER_9_194 VPWR VGND sg13g2_fill_1
X_08080_ _02221_ _02327_ _02346_ VPWR VGND sg13g2_nor2_1
XFILLER_115_711 VPWR VGND sg13g2_decap_4
XFILLER_54_0 VPWR VGND sg13g2_decap_8
XFILLER_114_221 VPWR VGND sg13g2_decap_8
XFILLER_115_788 VPWR VGND sg13g2_decap_8
X_08982_ VPWR _03168_ acc_sub.add_renorm0.exp\[0\] VGND sg13g2_inv_1
XFILLER_103_939 VPWR VGND sg13g2_decap_8
XFILLER_87_105 VPWR VGND sg13g2_decap_8
XFILLER_114_298 VPWR VGND sg13g2_decap_8
XFILLER_111_950 VPWR VGND sg13g2_decap_8
XFILLER_69_864 VPWR VGND sg13g2_decap_8
X_07933_ VPWR _02208_ fp16_sum_pipe.exp_mant_logic0.a\[9\] VGND sg13g2_inv_1
X_07864_ _02154_ _02155_ _02157_ _02158_ VPWR VGND sg13g2_nor3_1
XFILLER_96_672 VPWR VGND sg13g2_decap_8
XFILLER_68_374 VPWR VGND sg13g2_decap_8
XFILLER_3_91 VPWR VGND sg13g2_decap_8
X_09603_ VGND VPWR _03719_ _03696_ _03720_ _03694_ sg13g2_a21oi_1
X_07795_ _02094_ _01975_ net1747 VPWR VGND sg13g2_nand2_1
XFILLER_84_867 VPWR VGND sg13g2_fill_1
XFILLER_37_750 VPWR VGND sg13g2_decap_4
X_09534_ _03621_ acc_sum.add_renorm0.mantisa\[4\] _03651_ VPWR VGND sg13g2_nor2b_1
XFILLER_71_539 VPWR VGND sg13g2_fill_1
XFILLER_71_528 VPWR VGND sg13g2_decap_8
XFILLER_43_208 VPWR VGND sg13g2_fill_2
XFILLER_36_271 VPWR VGND sg13g2_fill_2
XFILLER_24_411 VPWR VGND sg13g2_decap_8
X_09465_ _03594_ VPWR _01253_ VGND net1915 _03593_ sg13g2_o21ai_1
XFILLER_19_1006 VPWR VGND sg13g2_decap_8
XFILLER_25_945 VPWR VGND sg13g2_decap_8
XFILLER_52_786 VPWR VGND sg13g2_fill_2
XFILLER_11_105 VPWR VGND sg13g2_decap_8
XFILLER_12_628 VPWR VGND sg13g2_decap_4
XFILLER_24_477 VPWR VGND sg13g2_decap_8
XFILLER_51_285 VPWR VGND sg13g2_decap_8
X_09396_ _01270_ _03538_ _03542_ VPWR VGND sg13g2_nand2_1
XFILLER_24_499 VPWR VGND sg13g2_decap_8
X_08278_ _02527_ _02526_ _02475_ VPWR VGND sg13g2_nand2_1
XFILLER_20_683 VPWR VGND sg13g2_decap_4
XFILLER_22_56 VPWR VGND sg13g2_decap_8
XFILLER_125_519 VPWR VGND sg13g2_fill_2
X_07229_ _01600_ _01599_ _01565_ VPWR VGND sg13g2_nand2_1
XFILLER_98_38 VPWR VGND sg13g2_decap_8
X_10240_ _04309_ _04310_ _04311_ _04312_ VPWR VGND sg13g2_nor3_1
XFILLER_79_639 VPWR VGND sg13g2_decap_4
X_10171_ _04248_ _04249_ _04250_ _04251_ VPWR VGND sg13g2_nor3_1
XFILLER_120_224 VPWR VGND sg13g2_decap_8
Xfanout140 net141 net140 VPWR VGND sg13g2_buf_2
XFILLER_59_330 VPWR VGND sg13g2_fill_1
XFILLER_102_972 VPWR VGND sg13g2_decap_8
X_13930_ VPWR _00481_ net7 VGND sg13g2_inv_1
XFILLER_74_311 VPWR VGND sg13g2_decap_8
XFILLER_19_227 VPWR VGND sg13g2_decap_8
XFILLER_90_804 VPWR VGND sg13g2_decap_8
XFILLER_75_889 VPWR VGND sg13g2_decap_8
XFILLER_47_75 VPWR VGND sg13g2_decap_8
X_13861_ VPWR _00412_ net47 VGND sg13g2_inv_1
X_12812_ acc\[13\] net1908 net1767 _06595_ VPWR VGND sg13g2_nand3_1
XFILLER_62_517 VPWR VGND sg13g2_fill_1
X_13792_ VPWR _00343_ net19 VGND sg13g2_inv_1
XFILLER_28_772 VPWR VGND sg13g2_fill_2
XFILLER_103_92 VPWR VGND sg13g2_decap_4
X_12743_ fpmul.reg_b_out\[14\] fp16_res_pipe.x2\[14\] net1952 _00924_ VPWR VGND sg13g2_mux2_1
XFILLER_42_230 VPWR VGND sg13g2_fill_1
XFILLER_16_945 VPWR VGND sg13g2_decap_8
XFILLER_43_786 VPWR VGND sg13g2_decap_8
XFILLER_43_764 VPWR VGND sg13g2_decap_8
XFILLER_15_455 VPWR VGND sg13g2_fill_1
XFILLER_15_477 VPWR VGND sg13g2_decap_8
X_12674_ _06487_ VPWR _00938_ VGND _06485_ net1741 sg13g2_o21ai_1
X_14413_ _00214_ VGND VPWR _00952_ fpmul.reg_a_out\[10\] clknet_leaf_127_clk sg13g2_dfrbpq_2
XFILLER_42_296 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
XFILLER_30_425 VPWR VGND sg13g2_fill_1
X_11625_ _05529_ VPWR _05530_ VGND fp16_sum_pipe.add_renorm0.mantisa\[11\] _05451_
+ sg13g2_o21ai_1
XFILLER_30_458 VPWR VGND sg13g2_fill_2
X_14344_ _00145_ VGND VPWR _00886_ fpmul.reg_p_out\[8\] clknet_leaf_88_clk sg13g2_dfrbpq_1
X_11556_ VPWR _05461_ _05459_ VGND sg13g2_inv_1
X_14275_ _00076_ VGND VPWR _00826_ fp16_res_pipe.x2\[8\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_10507_ _04550_ net1670 _04512_ VPWR VGND sg13g2_nand2_1
XFILLER_10_171 VPWR VGND sg13g2_decap_8
X_11487_ _05396_ VPWR _01033_ VGND net1945 _01766_ sg13g2_o21ai_1
X_13226_ _06951_ VPWR _00850_ VGND sipo.bit_counter\[0\] _06903_ sg13g2_o21ai_1
XFILLER_6_175 VPWR VGND sg13g2_decap_8
XFILLER_124_552 VPWR VGND sg13g2_fill_2
XFILLER_124_541 VPWR VGND sg13g2_decap_8
X_10438_ _04487_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[5\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[5\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_97_425 VPWR VGND sg13g2_fill_2
XFILLER_69_116 VPWR VGND sg13g2_fill_1
X_13157_ _06903_ _06880_ sipo.receiving VPWR VGND sg13g2_nand2_2
XFILLER_3_882 VPWR VGND sg13g2_decap_8
X_10369_ VPWR _04419_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[2\] VGND sg13g2_inv_1
XFILLER_100_909 VPWR VGND sg13g2_decap_8
XFILLER_85_609 VPWR VGND sg13g2_decap_8
XFILLER_69_138 VPWR VGND sg13g2_fill_1
X_13088_ _06850_ VPWR _00887_ VGND net1861 _06644_ sg13g2_o21ai_1
X_12108_ VPWR _05954_ _05953_ VGND sg13g2_inv_1
XFILLER_2_381 VPWR VGND sg13g2_decap_8
XFILLER_111_268 VPWR VGND sg13g2_fill_1
XFILLER_97_469 VPWR VGND sg13g2_decap_4
XFILLER_84_108 VPWR VGND sg13g2_decap_8
X_12039_ _05885_ net1857 net1864 VPWR VGND sg13g2_nand2_1
XFILLER_66_845 VPWR VGND sg13g2_fill_1
XFILLER_65_300 VPWR VGND sg13g2_decap_4
XFILLER_65_333 VPWR VGND sg13g2_fill_1
Xclkbuf_4_1_0_clk clknet_0_clk clknet_4_1_0_clk VPWR VGND sg13g2_buf_8
XFILLER_26_709 VPWR VGND sg13g2_decap_8
X_07580_ _01894_ _01890_ net1687 VPWR VGND sg13g2_nand2_1
XFILLER_19_783 VPWR VGND sg13g2_fill_1
XFILLER_33_230 VPWR VGND sg13g2_fill_2
X_09250_ fp16_res_pipe.op_sign_logic0.mantisa_a\[2\] _03403_ _03404_ VPWR VGND sg13g2_nor2_1
XFILLER_22_926 VPWR VGND sg13g2_decap_8
X_08201_ VPWR _02457_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[10\] VGND sg13g2_inv_1
X_09181_ _03344_ acc_sub.x2\[7\] net1896 VPWR VGND sg13g2_nand2_1
XFILLER_21_447 VPWR VGND sg13g2_fill_2
XFILLER_119_335 VPWR VGND sg13g2_fill_2
X_08132_ _02261_ net1648 _02393_ VPWR VGND sg13g2_nor2_1
X_08063_ _02329_ _02328_ _02221_ VPWR VGND sg13g2_nand2_1
Xplace1810 acc_sum.exp_mant_logic0.a\[4\] net1810 VPWR VGND sg13g2_buf_2
Xplace1821 fp16_res_pipe.seg_reg1.q\[21\] net1821 VPWR VGND sg13g2_buf_2
Xplace1854 fpmul.reg_a_out\[6\] net1854 VPWR VGND sg13g2_buf_1
XFILLER_1_808 VPWR VGND sg13g2_decap_8
Xplace1832 fp16_res_pipe.reg2en.q\[0\] net1832 VPWR VGND sg13g2_buf_2
Xplace1843 fp16_sum_pipe.reg1en.q\[0\] net1843 VPWR VGND sg13g2_buf_1
XFILLER_103_703 VPWR VGND sg13g2_fill_1
XFILLER_88_425 VPWR VGND sg13g2_decap_4
Xplace1887 net1886 net1887 VPWR VGND sg13g2_buf_1
Xplace1865 fpmul.reg_b_out\[4\] net1865 VPWR VGND sg13g2_buf_2
Xplace1876 net1875 net1876 VPWR VGND sg13g2_buf_2
X_08965_ VPWR _03151_ _03150_ VGND sg13g2_inv_1
Xplace1898 net1897 net1898 VPWR VGND sg13g2_buf_2
XFILLER_124_14 VPWR VGND sg13g2_decap_8
XFILLER_97_970 VPWR VGND sg13g2_decap_8
XFILLER_76_609 VPWR VGND sg13g2_fill_1
XFILLER_75_108 VPWR VGND sg13g2_decap_4
X_07916_ _02185_ _02190_ _02191_ VPWR VGND sg13g2_nor2_1
X_08896_ _03083_ _02973_ _03006_ VPWR VGND sg13g2_nand2_1
XFILLER_112_1013 VPWR VGND sg13g2_fill_1
XFILLER_68_182 VPWR VGND sg13g2_decap_8
X_07847_ _02142_ _02018_ net1794 VPWR VGND sg13g2_nand2_1
XFILLER_29_569 VPWR VGND sg13g2_fill_2
X_07778_ net1640 VPWR _02079_ VGND _02074_ _02078_ sg13g2_o21ai_1
XFILLER_84_686 VPWR VGND sg13g2_decap_8
XFILLER_56_399 VPWR VGND sg13g2_decap_8
XFILLER_17_56 VPWR VGND sg13g2_decap_8
X_09517_ _03634_ acc_sum.add_renorm0.mantisa\[7\] VPWR VGND sg13g2_inv_2
XFILLER_72_859 VPWR VGND sg13g2_fill_2
XFILLER_25_753 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_decap_8
XFILLER_13_926 VPWR VGND sg13g2_decap_8
XFILLER_52_594 VPWR VGND sg13g2_decap_8
XFILLER_12_436 VPWR VGND sg13g2_fill_1
X_09448_ VPWR _03584_ fp16_res_pipe.add_renorm0.exp\[2\] VGND sg13g2_inv_1
XFILLER_40_778 VPWR VGND sg13g2_decap_8
XFILLER_40_767 VPWR VGND sg13g2_decap_4
XFILLER_8_418 VPWR VGND sg13g2_decap_8
X_09379_ _03527_ VPWR _01272_ VGND _03518_ _03525_ sg13g2_o21ai_1
XFILLER_12_469 VPWR VGND sg13g2_decap_8
XFILLER_33_77 VPWR VGND sg13g2_decap_8
X_11410_ _05351_ net1707 fpdiv.div_out\[3\] VPWR VGND sg13g2_nand2_1
X_12390_ net1860 fpmul.reg_b_out\[0\] _06228_ _06236_ VPWR VGND sg13g2_nand3_1
XFILLER_33_99 VPWR VGND sg13g2_decap_8
XFILLER_126_806 VPWR VGND sg13g2_decap_8
X_11341_ _05295_ _05294_ net1634 VPWR VGND sg13g2_nand2_1
XFILLER_119_891 VPWR VGND sg13g2_decap_8
X_14060_ VPWR _00611_ net80 VGND sg13g2_inv_1
X_11272_ _05234_ net1661 acc_sum.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_4_657 VPWR VGND sg13g2_decap_8
XFILLER_3_112 VPWR VGND sg13g2_decap_8
XFILLER_106_574 VPWR VGND sg13g2_fill_1
X_13011_ _06778_ VPWR _06779_ VGND _06750_ fpmul.seg_reg0.q\[9\] sg13g2_o21ai_1
X_10223_ _01197_ _04295_ _04296_ VPWR VGND sg13g2_nand2_1
XFILLER_3_189 VPWR VGND sg13g2_decap_8
X_10154_ _04235_ _04177_ fp16_res_pipe.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_88_981 VPWR VGND sg13g2_decap_8
XFILLER_0_863 VPWR VGND sg13g2_decap_8
X_14962_ _00763_ VGND VPWR _01482_ acc_sub.add_renorm0.mantisa\[6\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_2
XFILLER_59_182 VPWR VGND sg13g2_decap_8
XFILLER_48_834 VPWR VGND sg13g2_fill_2
X_10085_ _01209_ _04169_ _04170_ VPWR VGND sg13g2_nand2_1
X_14893_ _00694_ VGND VPWR _01413_ acc_sub.op_sign_logic0.mantisa_b\[3\] clknet_leaf_69_clk
+ sg13g2_dfrbpq_2
XFILLER_101_290 VPWR VGND sg13g2_decap_4
XFILLER_48_856 VPWR VGND sg13g2_decap_8
X_13913_ VPWR _00464_ net5 VGND sg13g2_inv_1
XFILLER_114_91 VPWR VGND sg13g2_decap_8
XFILLER_63_826 VPWR VGND sg13g2_decap_8
X_13844_ VPWR _00395_ net30 VGND sg13g2_inv_1
XFILLER_35_539 VPWR VGND sg13g2_fill_2
XFILLER_16_720 VPWR VGND sg13g2_fill_2
XFILLER_16_742 VPWR VGND sg13g2_decap_8
X_13775_ VPWR _00326_ net137 VGND sg13g2_inv_1
X_10987_ _04979_ VPWR _01116_ VGND net1926 _02194_ sg13g2_o21ai_1
XFILLER_95_7 VPWR VGND sg13g2_fill_1
X_12726_ _06530_ _06440_ _06531_ VPWR VGND sg13g2_xor2_1
XFILLER_15_274 VPWR VGND sg13g2_decap_8
XFILLER_16_797 VPWR VGND sg13g2_fill_2
XFILLER_90_72 VPWR VGND sg13g2_decap_8
X_12657_ _06410_ _06409_ _06473_ VPWR VGND sg13g2_and2_1
XFILLER_30_255 VPWR VGND sg13g2_fill_1
XFILLER_31_756 VPWR VGND sg13g2_decap_4
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_12_981 VPWR VGND sg13g2_decap_8
X_11608_ _05509_ _05510_ _05508_ _05513_ VPWR VGND _05512_ sg13g2_nand4_1
X_12588_ VPWR _06404_ _06403_ VGND sg13g2_inv_1
X_14327_ _00128_ VGND VPWR _00870_ sipo.word\[15\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_7_451 VPWR VGND sg13g2_fill_1
XFILLER_7_440 VPWR VGND sg13g2_decap_8
XFILLER_116_316 VPWR VGND sg13g2_decap_8
XFILLER_7_484 VPWR VGND sg13g2_decap_8
X_11539_ _05442_ _05444_ VPWR VGND sg13g2_inv_4
X_14258_ _00059_ VGND VPWR _00809_ acc_sub.x2\[7\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_125_872 VPWR VGND sg13g2_decap_8
XFILLER_112_511 VPWR VGND sg13g2_fill_2
XFILLER_112_500 VPWR VGND sg13g2_decap_8
X_14189_ VPWR _00740_ net104 VGND sg13g2_inv_1
X_13209_ _06940_ VPWR _00856_ VGND _06939_ net1714 sg13g2_o21ai_1
XFILLER_98_745 VPWR VGND sg13g2_decap_8
XFILLER_112_577 VPWR VGND sg13g2_decap_4
XFILLER_100_717 VPWR VGND sg13g2_fill_1
XFILLER_100_706 VPWR VGND sg13g2_decap_8
XFILLER_98_789 VPWR VGND sg13g2_decap_8
XFILLER_39_812 VPWR VGND sg13g2_decap_8
XFILLER_94_940 VPWR VGND sg13g2_decap_8
X_08750_ _02946_ VPWR _01320_ VGND net1898 _02945_ sg13g2_o21ai_1
X_07701_ _02008_ VPWR _02009_ VGND _01751_ _01979_ sg13g2_o21ai_1
X_08681_ VGND VPWR net1671 _02849_ _02897_ net1739 sg13g2_a21oi_1
XFILLER_66_642 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
X_07632_ _01946_ net1641 _01926_ VPWR VGND sg13g2_nand2b_1
XFILLER_65_174 VPWR VGND sg13g2_fill_1
XFILLER_65_152 VPWR VGND sg13g2_decap_8
XFILLER_39_889 VPWR VGND sg13g2_decap_8
XFILLER_53_347 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
X_07563_ VPWR _01877_ _01783_ VGND sg13g2_inv_1
XFILLER_41_509 VPWR VGND sg13g2_decap_8
X_09302_ _03456_ fp16_res_pipe.op_sign_logic0.s_b fp16_res_pipe.op_sign_logic0.add_sub
+ VPWR VGND sg13g2_xnor2_1
XFILLER_110_49 VPWR VGND sg13g2_decap_8
X_07494_ VPWR _01817_ _01816_ VGND sg13g2_inv_1
XFILLER_62_892 VPWR VGND sg13g2_decap_8
XFILLER_22_712 VPWR VGND sg13g2_decap_8
X_09233_ fp16_res_pipe.op_sign_logic0.mantisa_a\[6\] _03386_ _03387_ VPWR VGND sg13g2_nor2_2
X_09164_ _03332_ VPWR _01292_ VGND net1905 _03331_ sg13g2_o21ai_1
XFILLER_119_154 VPWR VGND sg13g2_decap_8
XFILLER_119_14 VPWR VGND sg13g2_decap_8
XFILLER_108_817 VPWR VGND sg13g2_decap_8
X_08115_ _02327_ _02320_ _02377_ VPWR VGND sg13g2_nor2_1
X_09095_ _03277_ _03209_ _03096_ _03278_ VPWR VGND sg13g2_a21o_1
X_08046_ _02312_ net1692 _02279_ VPWR VGND sg13g2_nand2_1
XFILLER_122_308 VPWR VGND sg13g2_fill_2
XFILLER_115_360 VPWR VGND sg13g2_decap_8
Xplace1640 _02063_ net1640 VPWR VGND sg13g2_buf_2
Xplace1651 _01923_ net1651 VPWR VGND sg13g2_buf_2
Xplace1662 _04105_ net1662 VPWR VGND sg13g2_buf_2
XFILLER_77_907 VPWR VGND sg13g2_decap_4
Xplace1695 net1693 net1695 VPWR VGND sg13g2_buf_2
XFILLER_0_126 VPWR VGND sg13g2_decap_8
Xplace1684 _02250_ net1684 VPWR VGND sg13g2_buf_2
Xplace1673 _04460_ net1673 VPWR VGND sg13g2_buf_2
XFILLER_95_39 VPWR VGND sg13g2_decap_4
XFILLER_89_767 VPWR VGND sg13g2_decap_8
XFILLER_88_266 VPWR VGND sg13g2_decap_8
X_09997_ VGND VPWR _04084_ _04007_ _04085_ _04006_ sg13g2_a21oi_1
X_08948_ _02965_ _03134_ _03135_ VPWR VGND sg13g2_nor2_2
XFILLER_76_439 VPWR VGND sg13g2_fill_2
XFILLER_48_119 VPWR VGND sg13g2_decap_8
X_08879_ _03066_ net1788 acc_sub.add_renorm0.mantisa\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_45_804 VPWR VGND sg13g2_decap_4
XFILLER_84_450 VPWR VGND sg13g2_decap_8
XFILLER_57_675 VPWR VGND sg13g2_fill_1
X_10910_ _04919_ _04915_ _04811_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_77 VPWR VGND sg13g2_decap_8
X_11890_ fpdiv.divider0.counter\[0\] net1718 _05776_ VPWR VGND sg13g2_nor2_1
XFILLER_72_645 VPWR VGND sg13g2_decap_4
XFILLER_72_634 VPWR VGND sg13g2_fill_1
XFILLER_71_100 VPWR VGND sg13g2_fill_2
XFILLER_56_196 VPWR VGND sg13g2_fill_2
XFILLER_17_539 VPWR VGND sg13g2_decap_4
XFILLER_44_21 VPWR VGND sg13g2_decap_8
X_10841_ _04785_ VPWR _04853_ VGND _04817_ _04852_ sg13g2_o21ai_1
X_13560_ VPWR _00111_ net21 VGND sg13g2_inv_1
X_10772_ VGND VPWR net1709 _04782_ _04784_ _04783_ sg13g2_a21oi_1
XFILLER_25_572 VPWR VGND sg13g2_fill_2
X_13491_ VPWR _00042_ net83 VGND sg13g2_inv_1
X_12511_ VGND VPWR _06339_ net1953 _00953_ _06340_ sg13g2_a21oi_1
XFILLER_44_98 VPWR VGND sg13g2_decap_8
X_12442_ _06288_ _06286_ _06287_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_266 VPWR VGND sg13g2_decap_8
XFILLER_12_277 VPWR VGND sg13g2_fill_1
XFILLER_121_0 VPWR VGND sg13g2_decap_8
XFILLER_100_93 VPWR VGND sg13g2_decap_8
XFILLER_60_53 VPWR VGND sg13g2_fill_1
X_12373_ _06217_ _06218_ _06219_ VPWR VGND sg13g2_nor2_1
X_11324_ _03351_ _05176_ _05279_ VPWR VGND sg13g2_nor2_1
XFILLER_5_955 VPWR VGND sg13g2_decap_8
X_14112_ VPWR _00663_ net44 VGND sg13g2_inv_1
XFILLER_125_168 VPWR VGND sg13g2_decap_8
XFILLER_107_872 VPWR VGND sg13g2_fill_1
X_14043_ VPWR _00594_ net81 VGND sg13g2_inv_1
XFILLER_79_200 VPWR VGND sg13g2_decap_8
X_11255_ _05219_ acc_sum.exp_mant_logic0.a\[0\] net1680 acc_sum.op_sign_logic0.mantisa_a\[3\]
+ net1759 VPWR VGND sg13g2_a22oi_1
XFILLER_4_476 VPWR VGND sg13g2_decap_8
XFILLER_106_382 VPWR VGND sg13g2_decap_8
XFILLER_79_211 VPWR VGND sg13g2_fill_1
X_10206_ _01199_ _04280_ _04281_ VPWR VGND sg13g2_nand2_1
XFILLER_122_875 VPWR VGND sg13g2_decap_8
XFILLER_95_704 VPWR VGND sg13g2_decap_8
XFILLER_79_244 VPWR VGND sg13g2_decap_8
X_11186_ _05155_ _05124_ net1808 VPWR VGND sg13g2_nand2_1
XFILLER_79_299 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
X_10137_ _04219_ _04213_ _04218_ VPWR VGND sg13g2_nand2_1
XFILLER_94_247 VPWR VGND sg13g2_decap_4
X_14945_ _00746_ VGND VPWR _01465_ acc_sub.exp_mant_logic0.a\[13\] clknet_leaf_55_clk
+ sg13g2_dfrbpq_1
XFILLER_76_962 VPWR VGND sg13g2_decap_8
XFILLER_10_7 VPWR VGND sg13g2_decap_8
X_10068_ _04155_ _04126_ net1827 VPWR VGND sg13g2_nand2_1
XFILLER_63_601 VPWR VGND sg13g2_decap_4
XFILLER_91_954 VPWR VGND sg13g2_decap_8
X_14876_ _00677_ VGND VPWR _01396_ acc_sub.exp_mant_logic0.b\[2\] clknet_leaf_57_clk
+ sg13g2_dfrbpq_2
XFILLER_75_494 VPWR VGND sg13g2_fill_2
XFILLER_75_483 VPWR VGND sg13g2_fill_1
XFILLER_63_678 VPWR VGND sg13g2_fill_1
XFILLER_62_144 VPWR VGND sg13g2_decap_8
X_13827_ VPWR _00378_ net10 VGND sg13g2_inv_1
XFILLER_90_497 VPWR VGND sg13g2_decap_4
X_13758_ VPWR _00309_ net108 VGND sg13g2_inv_1
XFILLER_62_199 VPWR VGND sg13g2_decap_4
X_12709_ VPWR _06516_ div_result\[5\] VGND sg13g2_inv_1
X_13689_ VPWR _00240_ net65 VGND sg13g2_inv_1
XFILLER_116_124 VPWR VGND sg13g2_decap_8
XFILLER_104_308 VPWR VGND sg13g2_decap_8
X_09920_ _04017_ _04011_ _04016_ VPWR VGND sg13g2_nand2_2
X_09851_ _03740_ _03960_ _03961_ VPWR VGND sg13g2_nor2_1
X_08802_ acc_sub.add_renorm0.mantisa\[9\] _02988_ _02984_ _02989_ VPWR VGND sg13g2_nand3_1
XFILLER_113_886 VPWR VGND sg13g2_decap_8
XFILLER_100_503 VPWR VGND sg13g2_fill_1
X_09782_ _03822_ _03819_ _03897_ VPWR VGND sg13g2_nor2_1
XFILLER_85_225 VPWR VGND sg13g2_decap_8
XFILLER_100_569 VPWR VGND sg13g2_decap_8
XFILLER_85_236 VPWR VGND sg13g2_decap_8
XFILLER_67_962 VPWR VGND sg13g2_decap_4
XFILLER_67_940 VPWR VGND sg13g2_fill_1
X_08733_ VPWR _02935_ acc_sum.exp_mant_logic0.a\[14\] VGND sg13g2_inv_1
XFILLER_66_472 VPWR VGND sg13g2_decap_8
X_08664_ net1818 acc_sum.add_renorm0.mantisa\[7\] _02883_ VPWR VGND sg13g2_nor2_1
XFILLER_94_792 VPWR VGND sg13g2_fill_1
XFILLER_82_954 VPWR VGND sg13g2_decap_8
X_07615_ _01929_ _01920_ _01928_ VPWR VGND sg13g2_nand2_1
X_08595_ VPWR _02818_ _02817_ VGND sg13g2_inv_1
X_07546_ _01861_ _01862_ _01860_ _01433_ VPWR VGND sg13g2_nand3_1
XFILLER_53_177 VPWR VGND sg13g2_fill_2
XFILLER_41_328 VPWR VGND sg13g2_decap_4
XFILLER_14_35 VPWR VGND sg13g2_decap_8
X_07477_ acc_sub.exp_mant_logic0.a\[11\] _01799_ _01800_ VPWR VGND sg13g2_nor2_1
X_09216_ VPWR _03370_ fp16_res_pipe.op_sign_logic0.mantisa_a\[8\] VGND sg13g2_inv_1
X_09147_ VGND VPWR _03054_ net1800 _01299_ _03322_ sg13g2_a21oi_1
X_09078_ _03187_ _03157_ _03179_ _03262_ VPWR VGND sg13g2_nor3_1
XFILLER_108_647 VPWR VGND sg13g2_decap_8
XFILLER_5_229 VPWR VGND sg13g2_decap_8
XFILLER_30_56 VPWR VGND sg13g2_decap_8
XFILLER_122_105 VPWR VGND sg13g2_decap_8
X_08029_ _02233_ net1692 _02295_ VPWR VGND sg13g2_nor2_1
XFILLER_2_947 VPWR VGND sg13g2_decap_8
X_11040_ acc_sum.exp_mant_logic0.b\[8\] acc_sum.exp_mant_logic0.a\[8\] _05019_ VPWR
+ VGND sg13g2_xor2_1
XFILLER_39_21 VPWR VGND sg13g2_decap_8
XFILLER_7_1007 VPWR VGND sg13g2_decap_8
XFILLER_1_457 VPWR VGND sg13g2_decap_8
XFILLER_76_236 VPWR VGND sg13g2_fill_1
XFILLER_58_940 VPWR VGND sg13g2_fill_1
XFILLER_39_98 VPWR VGND sg13g2_decap_8
X_12991_ VPWR _06759_ _06758_ VGND sg13g2_inv_1
XFILLER_57_461 VPWR VGND sg13g2_fill_2
XFILLER_18_804 VPWR VGND sg13g2_decap_8
XFILLER_29_141 VPWR VGND sg13g2_decap_8
XFILLER_91_239 VPWR VGND sg13g2_decap_8
XFILLER_73_932 VPWR VGND sg13g2_fill_2
XFILLER_55_42 VPWR VGND sg13g2_decap_8
XFILLER_45_623 VPWR VGND sg13g2_fill_1
X_11942_ VPWR _05805_ fpmul.seg_reg0.q\[32\] VGND sg13g2_inv_1
XFILLER_17_325 VPWR VGND sg13g2_decap_8
X_14730_ _00531_ VGND VPWR _01258_ fp16_res_pipe.add_renorm0.exp\[1\] clknet_5_2__leaf_clk
+ sg13g2_dfrbpq_2
XFILLER_73_987 VPWR VGND sg13g2_fill_1
XFILLER_45_678 VPWR VGND sg13g2_decap_8
X_11873_ add_result\[1\] _05555_ net1850 _01014_ VPWR VGND sg13g2_mux2_1
XFILLER_44_133 VPWR VGND sg13g2_decap_8
X_14661_ _00462_ VGND VPWR _01189_ fp16_res_pipe.exp_mant_logic0.b\[14\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
X_13612_ VPWR _00163_ net111 VGND sg13g2_inv_1
X_14592_ _00393_ VGND VPWR _01124_ fp16_res_pipe.y\[3\] clknet_leaf_128_clk sg13g2_dfrbpq_1
XFILLER_44_188 VPWR VGND sg13g2_decap_4
X_10824_ VPWR _04836_ _04835_ VGND sg13g2_inv_1
XFILLER_26_870 VPWR VGND sg13g2_fill_1
XFILLER_125_1012 VPWR VGND sg13g2_fill_2
XFILLER_111_70 VPWR VGND sg13g2_decap_8
X_13543_ VPWR _00094_ net97 VGND sg13g2_inv_1
XFILLER_13_520 VPWR VGND sg13g2_fill_2
XFILLER_13_531 VPWR VGND sg13g2_fill_1
XFILLER_40_361 VPWR VGND sg13g2_decap_8
X_10755_ _04767_ VPWR _04768_ VGND net1822 _04762_ sg13g2_o21ai_1
X_13474_ VPWR _00025_ net33 VGND sg13g2_inv_1
X_10686_ _04699_ _04670_ _04681_ VPWR VGND sg13g2_nand2_1
X_12425_ _06270_ VPWR _06271_ VGND fpmul.reg_a_out\[5\] _06254_ sg13g2_o21ai_1
XFILLER_127_967 VPWR VGND sg13g2_decap_8
XFILLER_126_444 VPWR VGND sg13g2_fill_2
X_12356_ _06202_ _06201_ _06198_ VPWR VGND sg13g2_nand2b_1
XFILLER_126_477 VPWR VGND sg13g2_fill_1
XFILLER_58_7 VPWR VGND sg13g2_decap_8
X_11307_ _05265_ net1812 net1681 acc_sum.op_sign_logic0.mantisa_b\[8\] net1762 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_4_251 VPWR VGND sg13g2_fill_1
XFILLER_113_105 VPWR VGND sg13g2_decap_8
X_12287_ _06126_ _06132_ _06124_ _06133_ VPWR VGND sg13g2_nand3_1
XFILLER_5_785 VPWR VGND sg13g2_decap_8
XFILLER_122_661 VPWR VGND sg13g2_fill_2
XFILLER_110_801 VPWR VGND sg13g2_decap_8
X_14026_ VPWR _00577_ net98 VGND sg13g2_inv_1
X_11238_ _01088_ _05201_ _05202_ VPWR VGND sg13g2_nand2_1
XFILLER_45_1013 VPWR VGND sg13g2_fill_1
XFILLER_122_672 VPWR VGND sg13g2_fill_2
XFILLER_95_523 VPWR VGND sg13g2_decap_8
Xclkbuf_5_27__f_clk clknet_4_13_0_clk clknet_5_27__leaf_clk VPWR VGND sg13g2_buf_8
X_11169_ _05124_ _05136_ _05138_ VPWR VGND sg13g2_nor2_1
XFILLER_121_182 VPWR VGND sg13g2_decap_8
XFILLER_110_878 VPWR VGND sg13g2_decap_8
XFILLER_49_995 VPWR VGND sg13g2_decap_8
X_14928_ _00729_ VGND VPWR _01448_ fpdiv.divider0.divisor_reg\[8\] clknet_leaf_85_clk
+ sg13g2_dfrbpq_2
XFILLER_75_280 VPWR VGND sg13g2_decap_4
X_14859_ _00660_ VGND VPWR _01383_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[10\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_1
X_07400_ _01742_ net1890 acc\[6\] VPWR VGND sg13g2_nand2_1
X_08380_ _02619_ _02564_ _07116_ VPWR VGND sg13g2_nor2b_1
XFILLER_51_637 VPWR VGND sg13g2_fill_1
XFILLER_35_188 VPWR VGND sg13g2_decap_8
XFILLER_17_870 VPWR VGND sg13g2_decap_8
X_07331_ _01693_ net1666 _01625_ VPWR VGND sg13g2_nand2_1
XFILLER_50_147 VPWR VGND sg13g2_decap_8
XFILLER_118_901 VPWR VGND sg13g2_decap_8
X_07262_ _01631_ VPWR _01632_ VGND _01530_ _01630_ sg13g2_o21ai_1
XFILLER_84_0 VPWR VGND sg13g2_decap_8
X_07193_ VPWR _01565_ _01564_ VGND sg13g2_inv_1
X_09001_ VGND VPWR _03186_ _03187_ _03185_ net1699 sg13g2_a21oi_2
XFILLER_118_978 VPWR VGND sg13g2_decap_8
XFILLER_117_488 VPWR VGND sg13g2_decap_8
XFILLER_6_91 VPWR VGND sg13g2_decap_8
XFILLER_116_26 VPWR VGND sg13g2_decap_8
XFILLER_99_873 VPWR VGND sg13g2_decap_8
X_09903_ VPWR _04000_ fp16_res_pipe.exp_mant_logic0.b\[13\] VGND sg13g2_inv_1
XFILLER_99_884 VPWR VGND sg13g2_fill_1
XFILLER_98_383 VPWR VGND sg13g2_decap_8
X_09834_ VPWR _03945_ acc_sum.y\[9\] VGND sg13g2_inv_1
XFILLER_86_512 VPWR VGND sg13g2_fill_2
XFILLER_59_748 VPWR VGND sg13g2_decap_8
XFILLER_58_203 VPWR VGND sg13g2_decap_8
XFILLER_101_856 VPWR VGND sg13g2_decap_8
X_09765_ _03881_ _03880_ _03858_ VPWR VGND sg13g2_nand2_1
X_09696_ _03811_ VPWR _03812_ VGND _02806_ _03810_ sg13g2_o21ai_1
X_08716_ _02925_ net1819 acc_sum.seg_reg0.q\[27\] VPWR VGND sg13g2_nand2_1
XFILLER_67_792 VPWR VGND sg13g2_fill_2
XFILLER_39_494 VPWR VGND sg13g2_decap_8
X_08647_ _02867_ VPWR _02868_ VGND _02863_ _02866_ sg13g2_o21ai_1
XFILLER_92_29 VPWR VGND sg13g2_decap_8
XFILLER_82_740 VPWR VGND sg13g2_decap_8
XFILLER_54_464 VPWR VGND sg13g2_decap_8
XFILLER_15_807 VPWR VGND sg13g2_fill_2
XFILLER_70_935 VPWR VGND sg13g2_decap_4
X_08578_ VPWR _02802_ acc_sum.op_sign_logic0.s_a VGND sg13g2_inv_1
XFILLER_25_56 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_fill_1
X_07529_ _01850_ _01847_ acc_sub.exp_mant_logic0.a\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_23_884 VPWR VGND sg13g2_decap_8
XFILLER_50_681 VPWR VGND sg13g2_fill_1
X_10540_ VGND VPWR _04577_ net1849 _01162_ _04578_ sg13g2_a21oi_1
XFILLER_108_411 VPWR VGND sg13g2_decap_8
XFILLER_6_516 VPWR VGND sg13g2_decap_8
X_10471_ _04496_ VPWR _04519_ VGND _04517_ _04518_ sg13g2_o21ai_1
XFILLER_109_956 VPWR VGND sg13g2_decap_8
X_12210_ _06056_ _06053_ _06055_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_77 VPWR VGND sg13g2_decap_8
XFILLER_108_466 VPWR VGND sg13g2_decap_8
X_13190_ _06928_ net1712 sipo.word\[7\] VPWR VGND sg13g2_nand2_1
X_12141_ _05987_ net1866 _05982_ VPWR VGND sg13g2_xnor2_1
XFILLER_111_609 VPWR VGND sg13g2_decap_4
X_12072_ _05915_ _05917_ _05914_ _05918_ VPWR VGND sg13g2_nand3_1
XFILLER_103_160 VPWR VGND sg13g2_decap_8
XFILLER_89_361 VPWR VGND sg13g2_decap_4
X_11023_ VPWR _05002_ _05001_ VGND sg13g2_inv_1
XFILLER_77_534 VPWR VGND sg13g2_fill_1
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_65_729 VPWR VGND sg13g2_decap_4
XFILLER_49_258 VPWR VGND sg13g2_decap_8
X_12974_ _06744_ _06743_ net1961 VPWR VGND sg13g2_nand2_1
XFILLER_66_74 VPWR VGND sg13g2_decap_8
XFILLER_46_943 VPWR VGND sg13g2_decap_8
XFILLER_46_965 VPWR VGND sg13g2_fill_1
X_11925_ _05794_ net1879 fpmul.reg_b_out\[14\] VPWR VGND sg13g2_nand2_1
X_14713_ _00514_ VGND VPWR _01241_ fp16_res_pipe.exp_mant_logic0.a\[0\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
XFILLER_17_155 VPWR VGND sg13g2_decap_4
XFILLER_122_91 VPWR VGND sg13g2_decap_8
XFILLER_61_935 VPWR VGND sg13g2_decap_4
XFILLER_82_62 VPWR VGND sg13g2_decap_8
X_11856_ _05753_ VPWR _01021_ VGND net1756 _05752_ sg13g2_o21ai_1
X_14644_ _00445_ VGND VPWR net1833 fp16_res_pipe.reg3en.q\[0\] clknet_leaf_130_clk
+ sg13g2_dfrbpq_2
XFILLER_60_489 VPWR VGND sg13g2_fill_1
XFILLER_60_478 VPWR VGND sg13g2_decap_8
X_11787_ _05683_ _05689_ _05690_ VPWR VGND sg13g2_and2_1
X_14575_ _00376_ VGND VPWR _01107_ fp16_sum_pipe.exp_mant_logic0.b\[2\] clknet_leaf_135_clk
+ sg13g2_dfrbpq_2
X_10807_ _04819_ _04813_ _04818_ VPWR VGND sg13g2_nand2_1
X_13526_ VPWR _00077_ net35 VGND sg13g2_inv_1
XFILLER_41_692 VPWR VGND sg13g2_fill_1
XFILLER_41_681 VPWR VGND sg13g2_decap_8
XFILLER_9_343 VPWR VGND sg13g2_decap_8
XFILLER_13_394 VPWR VGND sg13g2_decap_8
XFILLER_14_895 VPWR VGND sg13g2_decap_8
X_10738_ _04750_ _04635_ _04751_ VPWR VGND sg13g2_and2_1
X_13457_ _07108_ net1752 sipo.shift_reg\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_40_191 VPWR VGND sg13g2_fill_1
XFILLER_9_354 VPWR VGND sg13g2_fill_1
XFILLER_9_365 VPWR VGND sg13g2_decap_4
X_12408_ _06254_ net1854 fpmul.reg_b_out\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_9_387 VPWR VGND sg13g2_decap_8
XFILLER_9_398 VPWR VGND sg13g2_fill_1
XFILLER_127_764 VPWR VGND sg13g2_decap_8
XFILLER_126_252 VPWR VGND sg13g2_decap_8
X_13388_ VGND VPWR _07003_ net1695 _00807_ _07070_ sg13g2_a21oi_1
X_12339_ _06183_ _06184_ _06185_ VPWR VGND _06181_ sg13g2_nand3b_1
XFILLER_123_981 VPWR VGND sg13g2_decap_8
X_14009_ VPWR _00560_ net19 VGND sg13g2_inv_1
XFILLER_122_491 VPWR VGND sg13g2_decap_8
X_07880_ _02167_ net1885 acc_sub.x2\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_96_887 VPWR VGND sg13g2_fill_1
XFILLER_95_375 VPWR VGND sg13g2_fill_2
XFILLER_37_910 VPWR VGND sg13g2_decap_8
X_09550_ _03667_ _03659_ _03652_ _03633_ VPWR VGND sg13g2_and3_2
XFILLER_110_697 VPWR VGND sg13g2_fill_1
XFILLER_95_397 VPWR VGND sg13g2_fill_2
XFILLER_95_386 VPWR VGND sg13g2_fill_1
X_08501_ VPWR _02726_ _02724_ VGND sg13g2_inv_1
XFILLER_52_902 VPWR VGND sg13g2_fill_2
XFILLER_37_987 VPWR VGND sg13g2_decap_8
XFILLER_36_453 VPWR VGND sg13g2_decap_8
X_09481_ _03605_ net1827 VPWR VGND sg13g2_inv_2
X_08432_ VGND VPWR _01772_ fpdiv.divider0.remainder_reg\[5\] _02666_ _02665_ sg13g2_a21oi_1
XFILLER_51_401 VPWR VGND sg13g2_decap_8
XFILLER_23_103 VPWR VGND sg13g2_fill_1
XFILLER_24_604 VPWR VGND sg13g2_decap_4
XFILLER_63_294 VPWR VGND sg13g2_fill_2
X_08363_ VPWR _02606_ instr\[3\] VGND sg13g2_inv_1
X_07314_ _01677_ VPWR _01678_ VGND _01571_ net1667 sg13g2_o21ai_1
X_08294_ _02469_ _02340_ _02541_ VPWR VGND sg13g2_nor2_1
X_07245_ _01615_ _01614_ _01583_ _01616_ VPWR VGND sg13g2_a21o_1
XFILLER_11_14 VPWR VGND sg13g2_decap_8
XFILLER_127_14 VPWR VGND sg13g2_decap_8
X_07176_ VPWR _01548_ acc_sub.op_sign_logic0.mantisa_a\[1\] VGND sg13g2_inv_1
XFILLER_118_775 VPWR VGND sg13g2_decap_8
XFILLER_117_252 VPWR VGND sg13g2_decap_8
XFILLER_106_915 VPWR VGND sg13g2_decap_8
XFILLER_105_436 VPWR VGND sg13g2_fill_2
XFILLER_120_439 VPWR VGND sg13g2_decap_4
XFILLER_113_480 VPWR VGND sg13g2_fill_2
XFILLER_101_653 VPWR VGND sg13g2_decap_8
X_09817_ VPWR _03930_ _03818_ VGND sg13g2_inv_1
XFILLER_100_152 VPWR VGND sg13g2_decap_4
XFILLER_86_364 VPWR VGND sg13g2_decap_4
XFILLER_19_409 VPWR VGND sg13g2_decap_8
Xclkbuf_5_10__f_clk clknet_4_5_0_clk clknet_5_10__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_28_910 VPWR VGND sg13g2_decap_8
XFILLER_100_174 VPWR VGND sg13g2_decap_8
X_09748_ _03863_ VPWR _03864_ VGND _02920_ net1690 sg13g2_o21ai_1
XFILLER_86_386 VPWR VGND sg13g2_fill_2
XFILLER_74_526 VPWR VGND sg13g2_decap_8
XFILLER_46_239 VPWR VGND sg13g2_decap_8
XFILLER_39_291 VPWR VGND sg13g2_decap_8
X_09679_ VGND VPWR _03793_ net1807 _03795_ _03794_ sg13g2_a21oi_1
XFILLER_82_570 VPWR VGND sg13g2_fill_2
XFILLER_70_710 VPWR VGND sg13g2_fill_2
XFILLER_61_209 VPWR VGND sg13g2_fill_2
XFILLER_54_250 VPWR VGND sg13g2_decap_8
XFILLER_36_77 VPWR VGND sg13g2_decap_8
X_11710_ _05614_ _05587_ _05613_ VPWR VGND sg13g2_xnor2_1
XFILLER_15_604 VPWR VGND sg13g2_fill_2
XFILLER_28_987 VPWR VGND sg13g2_decap_8
X_12690_ _06460_ _06420_ _06500_ VPWR VGND sg13g2_xor2_1
XFILLER_52_21 VPWR VGND sg13g2_decap_8
X_11641_ _05544_ _05545_ _05543_ _05546_ VPWR VGND sg13g2_nand3_1
X_14360_ _00161_ VGND VPWR _00902_ _00013_ clknet_leaf_87_clk sg13g2_dfrbpq_1
X_11572_ _05427_ _05476_ _05477_ VPWR VGND sg13g2_nor2_2
X_13311_ VGND VPWR net1677 _07020_ _00835_ _07021_ sg13g2_a21oi_1
XFILLER_7_825 VPWR VGND sg13g2_decap_8
X_10523_ net1673 VPWR _04564_ VGND _04420_ _04563_ sg13g2_o21ai_1
XFILLER_11_854 VPWR VGND sg13g2_decap_8
XFILLER_22_191 VPWR VGND sg13g2_decap_4
X_14291_ _00092_ VGND VPWR _00835_ acc\[1\] clknet_leaf_50_clk sg13g2_dfrbpq_2
X_13242_ _06967_ net1742 sipo.word\[15\] VPWR VGND sg13g2_nand2_1
X_10454_ _04474_ _04501_ _04429_ _04502_ VPWR VGND sg13g2_nor3_1
X_13173_ VPWR _06916_ sipo.shift_reg\[13\] VGND sg13g2_inv_1
X_10385_ VPWR _04435_ _04434_ VGND sg13g2_inv_1
XFILLER_124_767 VPWR VGND sg13g2_decap_8
X_12124_ _05968_ _05969_ _05970_ VPWR VGND sg13g2_nor2_1
XFILLER_123_266 VPWR VGND sg13g2_decap_8
XFILLER_112_929 VPWR VGND sg13g2_decap_8
XFILLER_2_563 VPWR VGND sg13g2_fill_2
XFILLER_117_91 VPWR VGND sg13g2_decap_8
XFILLER_78_854 VPWR VGND sg13g2_decap_8
XFILLER_77_40 VPWR VGND sg13g2_fill_1
X_12055_ _05901_ net1855 net1866 VPWR VGND sg13g2_nand2_1
XFILLER_78_887 VPWR VGND sg13g2_fill_2
XFILLER_38_718 VPWR VGND sg13g2_fill_1
X_11006_ _04989_ fp16_res_pipe.x2\[1\] net1925 VPWR VGND sg13g2_nand2_1
XFILLER_120_995 VPWR VGND sg13g2_decap_8
XFILLER_65_548 VPWR VGND sg13g2_decap_8
XFILLER_37_239 VPWR VGND sg13g2_decap_8
XFILLER_19_943 VPWR VGND sg13g2_decap_8
XFILLER_18_442 VPWR VGND sg13g2_fill_2
X_12957_ acc\[1\] load_en _03983_ _06728_ VPWR VGND sg13g2_nand3_1
XFILLER_45_272 VPWR VGND sg13g2_decap_8
XFILLER_18_486 VPWR VGND sg13g2_fill_1
X_12888_ _06665_ _06661_ _06664_ _06502_ net1949 VPWR VGND sg13g2_a22oi_1
XFILLER_61_732 VPWR VGND sg13g2_decap_4
X_11908_ VGND VPWR net1880 _05781_ _00998_ _05782_ sg13g2_a21oi_1
XFILLER_45_294 VPWR VGND sg13g2_decap_8
XFILLER_34_968 VPWR VGND sg13g2_decap_8
XFILLER_33_423 VPWR VGND sg13g2_fill_1
X_14627_ _00428_ VGND VPWR _01159_ fp16_sum_pipe.add_renorm0.exp\[6\] clknet_leaf_98_clk
+ sg13g2_dfrbpq_2
XFILLER_21_629 VPWR VGND sg13g2_decap_8
X_11839_ _05666_ _05662_ _05738_ VPWR VGND sg13g2_and2_1
XFILLER_33_478 VPWR VGND sg13g2_decap_8
XFILLER_20_106 VPWR VGND sg13g2_decap_8
X_14558_ _00359_ VGND VPWR _01094_ acc_sum.op_sign_logic0.mantisa_a\[10\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_9_140 VPWR VGND sg13g2_decap_8
X_13509_ VPWR _00060_ net34 VGND sg13g2_inv_1
X_14489_ _00290_ VGND VPWR _01027_ add_result\[14\] clknet_leaf_97_clk sg13g2_dfrbpq_2
XFILLER_127_583 VPWR VGND sg13g2_decap_8
XFILLER_114_200 VPWR VGND sg13g2_decap_8
XFILLER_115_767 VPWR VGND sg13g2_decap_8
X_08981_ _03167_ _03166_ _03163_ VPWR VGND sg13g2_nand2_1
XFILLER_114_277 VPWR VGND sg13g2_decap_8
XFILLER_69_810 VPWR VGND sg13g2_fill_2
XFILLER_87_139 VPWR VGND sg13g2_decap_8
XFILLER_69_854 VPWR VGND sg13g2_fill_1
XFILLER_69_843 VPWR VGND sg13g2_decap_8
X_07932_ _02204_ _02206_ _02207_ VPWR VGND sg13g2_nor2_1
X_07863_ _02156_ _02024_ _02157_ VPWR VGND sg13g2_nor2_1
XFILLER_84_813 VPWR VGND sg13g2_fill_1
XFILLER_68_353 VPWR VGND sg13g2_decap_8
XFILLER_56_504 VPWR VGND sg13g2_decap_8
XFILLER_3_70 VPWR VGND sg13g2_decap_8
XFILLER_29_718 VPWR VGND sg13g2_decap_8
X_09602_ _03692_ _03717_ _03719_ VPWR VGND sg13g2_nor2_1
XFILLER_95_161 VPWR VGND sg13g2_decap_8
XFILLER_84_824 VPWR VGND sg13g2_decap_8
XFILLER_56_537 VPWR VGND sg13g2_decap_8
XFILLER_56_515 VPWR VGND sg13g2_fill_1
XFILLER_28_239 VPWR VGND sg13g2_decap_8
XFILLER_113_49 VPWR VGND sg13g2_decap_8
X_09533_ VPWR _03650_ acc_sum.add_renorm0.mantisa\[5\] VGND sg13g2_inv_1
X_07794_ _02088_ _02090_ _02092_ _02093_ VPWR VGND sg13g2_nor3_1
XFILLER_56_559 VPWR VGND sg13g2_fill_1
XFILLER_58_1012 VPWR VGND sg13g2_fill_2
XFILLER_52_710 VPWR VGND sg13g2_fill_2
XFILLER_36_261 VPWR VGND sg13g2_fill_2
XFILLER_25_924 VPWR VGND sg13g2_decap_8
XFILLER_52_754 VPWR VGND sg13g2_decap_8
X_09464_ _03594_ acc_sub.x2\[12\] net1913 VPWR VGND sg13g2_nand2_1
X_08415_ _02643_ _02648_ _02650_ VPWR VGND sg13g2_nor2_2
XFILLER_51_264 VPWR VGND sg13g2_decap_8
X_09395_ VGND VPWR net1770 fp16_res_pipe.add_renorm0.mantisa\[5\] _03542_ _03541_
+ sg13g2_a21oi_1
X_08346_ _02588_ VPWR _02589_ VGND sipo.word_ready _02581_ sg13g2_o21ai_1
XFILLER_40_938 VPWR VGND sg13g2_decap_4
XFILLER_125_7 VPWR VGND sg13g2_decap_8
X_08277_ _02524_ _02525_ _02521_ _02526_ VPWR VGND sg13g2_nand3_1
XFILLER_22_35 VPWR VGND sg13g2_decap_8
X_07228_ _01598_ VPWR _01599_ VGND _01548_ _01550_ sg13g2_o21ai_1
X_07159_ VPWR _01531_ acc_sub.op_sign_logic0.mantisa_a\[5\] VGND sg13g2_inv_1
XFILLER_4_839 VPWR VGND sg13g2_decap_8
XFILLER_120_203 VPWR VGND sg13g2_decap_8
X_10170_ _03615_ _04233_ _04250_ VPWR VGND sg13g2_nor2_1
Xfanout130 net131 net130 VPWR VGND sg13g2_buf_1
XFILLER_102_951 VPWR VGND sg13g2_decap_8
XFILLER_93_109 VPWR VGND sg13g2_decap_4
Xfanout141 net2 net141 VPWR VGND sg13g2_buf_2
XFILLER_75_846 VPWR VGND sg13g2_fill_1
XFILLER_47_54 VPWR VGND sg13g2_decap_8
XFILLER_74_356 VPWR VGND sg13g2_decap_8
XFILLER_62_507 VPWR VGND sg13g2_decap_4
XFILLER_47_559 VPWR VGND sg13g2_decap_8
X_13860_ VPWR _00411_ net43 VGND sg13g2_inv_1
X_12811_ VGND VPWR net1935 add_result\[13\] _06594_ net1943 sg13g2_a21oi_1
X_13791_ VPWR _00342_ net20 VGND sg13g2_inv_1
XFILLER_16_924 VPWR VGND sg13g2_decap_8
XFILLER_27_250 VPWR VGND sg13g2_fill_2
XFILLER_83_890 VPWR VGND sg13g2_decap_8
X_12742_ fpmul.reg_b_out\[15\] fp16_res_pipe.x2\[15\] net1951 _00925_ VPWR VGND sg13g2_mux2_1
XFILLER_43_743 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_fill_2
XFILLER_27_283 VPWR VGND sg13g2_decap_8
X_12673_ _06479_ VPWR _06487_ VGND net1735 _06486_ sg13g2_o21ai_1
XFILLER_70_551 VPWR VGND sg13g2_decap_4
XFILLER_30_404 VPWR VGND sg13g2_decap_8
XFILLER_70_595 VPWR VGND sg13g2_decap_8
X_14412_ _00213_ VGND VPWR _00951_ fpmul.reg_a_out\[9\] clknet_leaf_92_clk sg13g2_dfrbpq_2
X_11624_ _05529_ fp16_sum_pipe.add_renorm0.mantisa\[11\] fp16_sum_pipe.add_renorm0.mantisa\[10\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_949 VPWR VGND sg13g2_decap_8
X_14343_ _00144_ VGND VPWR _00885_ fpmul.reg_p_out\[7\] clknet_leaf_81_clk sg13g2_dfrbpq_1
X_11486_ _05396_ fp16_res_pipe.x2\[4\] net1945 VPWR VGND sg13g2_nand2_1
X_14274_ _00075_ VGND VPWR _00825_ fp16_res_pipe.x2\[7\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_10506_ VGND VPWR _04548_ net1848 _01167_ _04549_ sg13g2_a21oi_1
XFILLER_109_594 VPWR VGND sg13g2_fill_1
XFILLER_109_583 VPWR VGND sg13g2_fill_2
XFILLER_109_572 VPWR VGND sg13g2_decap_8
XFILLER_109_561 VPWR VGND sg13g2_fill_1
X_13225_ _06951_ sipo.bit_counter\[0\] net3 VPWR VGND sg13g2_nand2_1
XFILLER_6_154 VPWR VGND sg13g2_decap_8
X_10437_ VGND VPWR _04483_ _04437_ _04486_ _04485_ sg13g2_a21oi_1
XFILLER_98_905 VPWR VGND sg13g2_decap_8
XFILLER_111_203 VPWR VGND sg13g2_fill_2
XFILLER_97_404 VPWR VGND sg13g2_decap_8
XFILLER_88_50 VPWR VGND sg13g2_decap_8
X_13156_ _06902_ _06901_ VPWR VGND sg13g2_inv_2
XFILLER_40_7 VPWR VGND sg13g2_decap_8
XFILLER_3_861 VPWR VGND sg13g2_decap_8
X_10368_ VGND VPWR _04412_ _04414_ _04418_ _04417_ sg13g2_a21oi_1
XFILLER_97_448 VPWR VGND sg13g2_fill_2
X_13087_ net1700 _06849_ _06809_ _06850_ VPWR VGND sg13g2_nand3_1
X_12107_ _05953_ net1860 fpmul.reg_b_out\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_2_360 VPWR VGND sg13g2_decap_8
X_10299_ _04367_ _04366_ net1636 VPWR VGND sg13g2_nand2_1
XFILLER_111_247 VPWR VGND sg13g2_decap_8
X_12038_ _05884_ _05882_ _05883_ VPWR VGND sg13g2_nand2_1
XFILLER_120_792 VPWR VGND sg13g2_decap_8
XFILLER_93_610 VPWR VGND sg13g2_decap_4
XFILLER_77_183 VPWR VGND sg13g2_decap_8
XFILLER_38_537 VPWR VGND sg13g2_decap_8
XFILLER_92_175 VPWR VGND sg13g2_decap_4
XFILLER_80_315 VPWR VGND sg13g2_fill_1
X_13989_ VPWR _00540_ net9 VGND sg13g2_inv_1
XFILLER_92_197 VPWR VGND sg13g2_decap_8
XFILLER_61_551 VPWR VGND sg13g2_fill_2
XFILLER_61_540 VPWR VGND sg13g2_decap_8
XFILLER_21_404 VPWR VGND sg13g2_decap_8
XFILLER_22_905 VPWR VGND sg13g2_decap_8
XFILLER_61_595 VPWR VGND sg13g2_decap_8
X_08200_ _01373_ _02455_ _02456_ VPWR VGND sg13g2_nand2_1
XFILLER_21_415 VPWR VGND sg13g2_fill_2
X_09180_ _03343_ acc_sum.exp_mant_logic0.b\[7\] VPWR VGND sg13g2_inv_2
XFILLER_119_314 VPWR VGND sg13g2_decap_8
X_08131_ _02269_ net1652 _02392_ VPWR VGND sg13g2_nor2_1
X_08062_ VPWR _02328_ _02327_ VGND sg13g2_inv_1
Xplace1800 acc_sub.reg3en.q\[0\] net1800 VPWR VGND sg13g2_buf_1
Xplace1811 acc_sum.exp_mant_logic0.b\[6\] net1811 VPWR VGND sg13g2_buf_2
Xplace1822 fp16_res_pipe.seg_reg1.q\[21\] net1822 VPWR VGND sg13g2_buf_2
Xplace1844 fp16_sum_pipe.reg2en.q\[0\] net1844 VPWR VGND sg13g2_buf_1
Xplace1833 net1832 net1833 VPWR VGND sg13g2_buf_2
XFILLER_115_586 VPWR VGND sg13g2_decap_8
XFILLER_103_726 VPWR VGND sg13g2_fill_1
XFILLER_89_916 VPWR VGND sg13g2_fill_1
XFILLER_88_404 VPWR VGND sg13g2_decap_8
Xplace1888 net1887 net1888 VPWR VGND sg13g2_buf_2
Xplace1855 fpmul.reg_a_out\[5\] net1855 VPWR VGND sg13g2_buf_2
Xplace1877 net1875 net1877 VPWR VGND sg13g2_buf_2
Xplace1866 fpmul.reg_b_out\[3\] net1866 VPWR VGND sg13g2_buf_2
X_08964_ _03150_ _01711_ _03142_ VPWR VGND sg13g2_xnor2_1
Xplace1899 net1898 net1899 VPWR VGND sg13g2_buf_2
XFILLER_102_269 VPWR VGND sg13g2_decap_8
XFILLER_102_247 VPWR VGND sg13g2_fill_2
X_07915_ _02190_ _02188_ _02189_ VPWR VGND sg13g2_nand2_1
X_08895_ _03006_ _02971_ _03082_ VPWR VGND sg13g2_nor2_1
XFILLER_84_621 VPWR VGND sg13g2_decap_8
XFILLER_68_161 VPWR VGND sg13g2_decap_8
X_07846_ _02089_ _01977_ _02141_ VPWR VGND sg13g2_nor2_1
XFILLER_83_131 VPWR VGND sg13g2_fill_2
XFILLER_29_548 VPWR VGND sg13g2_decap_8
X_07777_ _02076_ _02077_ _02075_ _02078_ VPWR VGND sg13g2_nand3_1
XFILLER_95_1009 VPWR VGND sg13g2_decap_4
XFILLER_72_827 VPWR VGND sg13g2_decap_8
XFILLER_16_209 VPWR VGND sg13g2_fill_2
XFILLER_17_35 VPWR VGND sg13g2_decap_8
X_09516_ _03633_ _03631_ VPWR VGND sg13g2_inv_2
XFILLER_72_849 VPWR VGND sg13g2_fill_2
XFILLER_13_905 VPWR VGND sg13g2_decap_8
X_09447_ _03583_ VPWR _01260_ VGND net1832 _03582_ sg13g2_o21ai_1
XFILLER_80_882 VPWR VGND sg13g2_decap_8
XFILLER_40_713 VPWR VGND sg13g2_decap_8
X_09378_ _03527_ net1738 _03526_ fp16_res_pipe.add_renorm0.mantisa\[7\] net1770 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_33_56 VPWR VGND sg13g2_decap_8
X_08329_ VPWR _02574_ _02573_ VGND sg13g2_inv_1
X_11340_ _05292_ _05293_ _05291_ _05294_ VPWR VGND sg13g2_nand3_1
XFILLER_119_870 VPWR VGND sg13g2_decap_8
X_13010_ _06778_ _06750_ fpmul.seg_reg0.q\[8\] VPWR VGND sg13g2_nand2b_1
X_11271_ _05233_ net1655 acc_sum.exp_mant_logic0.a\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_3_168 VPWR VGND sg13g2_decap_8
X_10222_ _04296_ fp16_res_pipe.exp_mant_logic0.b\[3\] net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[6\]
+ net1763 VPWR VGND sg13g2_a22oi_1
XFILLER_106_586 VPWR VGND sg13g2_decap_8
Xclkbuf_5_8__f_clk clknet_4_4_0_clk clknet_5_8__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_121_578 VPWR VGND sg13g2_fill_2
XFILLER_94_418 VPWR VGND sg13g2_fill_1
XFILLER_94_407 VPWR VGND sg13g2_decap_8
XFILLER_88_960 VPWR VGND sg13g2_decap_8
XFILLER_0_842 VPWR VGND sg13g2_decap_8
X_14961_ _00762_ VGND VPWR _01481_ acc_sub.add_renorm0.mantisa\[5\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_2
XFILLER_102_770 VPWR VGND sg13g2_decap_8
X_10084_ _04170_ fp16_res_pipe.exp_mant_logic0.a\[4\] net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[7\]
+ net1764 VPWR VGND sg13g2_a22oi_1
X_14892_ _00693_ VGND VPWR _01412_ acc_sub.op_sign_logic0.mantisa_b\[2\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_2
XFILLER_114_70 VPWR VGND sg13g2_decap_8
XFILLER_87_492 VPWR VGND sg13g2_decap_8
X_13912_ VPWR _00463_ net27 VGND sg13g2_inv_1
XFILLER_74_30 VPWR VGND sg13g2_decap_8
XFILLER_62_315 VPWR VGND sg13g2_decap_8
X_13843_ VPWR _00394_ net36 VGND sg13g2_inv_1
XFILLER_35_518 VPWR VGND sg13g2_decap_8
XFILLER_74_74 VPWR VGND sg13g2_decap_8
XFILLER_56_890 VPWR VGND sg13g2_decap_4
X_13774_ VPWR _00325_ net108 VGND sg13g2_inv_1
X_10986_ _04979_ fp16_res_pipe.x2\[11\] net1924 VPWR VGND sg13g2_nand2_1
XFILLER_15_231 VPWR VGND sg13g2_fill_1
XFILLER_16_776 VPWR VGND sg13g2_decap_8
X_12725_ _06530_ _06529_ _06447_ VPWR VGND sg13g2_nand2_1
XFILLER_43_595 VPWR VGND sg13g2_fill_2
XFILLER_30_212 VPWR VGND sg13g2_decap_8
XFILLER_88_7 VPWR VGND sg13g2_decap_4
X_12656_ _06471_ _06470_ _06472_ VPWR VGND sg13g2_xor2_1
XFILLER_31_746 VPWR VGND sg13g2_decap_4
X_12587_ _06397_ _06402_ _06403_ VPWR VGND sg13g2_nor2_1
XFILLER_12_960 VPWR VGND sg13g2_decap_8
X_11607_ VGND VPWR _05475_ _05428_ _05512_ _05511_ sg13g2_a21oi_1
XFILLER_30_267 VPWR VGND sg13g2_fill_2
X_14326_ _00127_ VGND VPWR _00869_ sipo.word\[14\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_11_481 VPWR VGND sg13g2_decap_8
XFILLER_116_328 VPWR VGND sg13g2_decap_8
XFILLER_116_306 VPWR VGND sg13g2_fill_1
XFILLER_8_986 VPWR VGND sg13g2_decap_8
XFILLER_7_463 VPWR VGND sg13g2_decap_8
XFILLER_125_851 VPWR VGND sg13g2_decap_8
XFILLER_99_60 VPWR VGND sg13g2_decap_8
X_11469_ fpdiv.reg_b_out\[12\] fp16_res_pipe.x2\[12\] net1939 _01041_ VPWR VGND sg13g2_mux2_1
X_14257_ _00058_ VGND VPWR _00808_ acc_sub.x2\[6\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_14188_ VPWR _00739_ net116 VGND sg13g2_inv_1
X_13208_ _06940_ net1714 sipo.word\[1\] VPWR VGND sg13g2_nand2_1
X_13139_ VPWR _06890_ _06889_ VGND sg13g2_inv_1
XFILLER_112_556 VPWR VGND sg13g2_decap_4
XFILLER_98_768 VPWR VGND sg13g2_decap_8
X_07700_ _02008_ _01959_ acc_sub.exp_mant_logic0.a\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_85_429 VPWR VGND sg13g2_decap_8
XFILLER_66_610 VPWR VGND sg13g2_decap_8
X_08680_ _02896_ net1668 _02769_ VPWR VGND sg13g2_nand2_1
XFILLER_65_131 VPWR VGND sg13g2_decap_8
XFILLER_39_868 VPWR VGND sg13g2_decap_8
XFILLER_38_345 VPWR VGND sg13g2_decap_8
XFILLER_94_996 VPWR VGND sg13g2_decap_8
XFILLER_93_462 VPWR VGND sg13g2_fill_1
XFILLER_81_602 VPWR VGND sg13g2_decap_4
X_07562_ VGND VPWR _01875_ _01834_ _01876_ _01794_ sg13g2_a21oi_1
XFILLER_80_112 VPWR VGND sg13g2_decap_8
XFILLER_19_570 VPWR VGND sg13g2_decap_4
XFILLER_110_28 VPWR VGND sg13g2_decap_8
X_07493_ _01814_ _01815_ _01816_ VPWR VGND sg13g2_nor2_1
XFILLER_80_189 VPWR VGND sg13g2_fill_1
XFILLER_80_178 VPWR VGND sg13g2_decap_8
X_09232_ VPWR _03386_ fp16_res_pipe.op_sign_logic0.mantisa_b\[6\] VGND sg13g2_inv_1
XFILLER_10_919 VPWR VGND sg13g2_decap_8
XFILLER_21_223 VPWR VGND sg13g2_fill_2
X_09163_ _03332_ acc_sub.x2\[13\] net1903 VPWR VGND sg13g2_nand2_1
XFILLER_119_133 VPWR VGND sg13g2_decap_8
XFILLER_9_91 VPWR VGND sg13g2_decap_8
X_08114_ _02268_ net1652 _02376_ VPWR VGND sg13g2_nor2_1
X_09094_ _03277_ _03207_ _03187_ VPWR VGND sg13g2_nand2_1
X_08045_ _02311_ _02207_ _02310_ VPWR VGND sg13g2_xnor2_1
XFILLER_116_884 VPWR VGND sg13g2_decap_8
Xplace1641 _01944_ net1641 VPWR VGND sg13g2_buf_2
Xplace1663 _05106_ net1663 VPWR VGND sg13g2_buf_2
Xplace1652 _02322_ net1652 VPWR VGND sg13g2_buf_1
XFILLER_115_394 VPWR VGND sg13g2_fill_1
Xplace1685 _01871_ net1685 VPWR VGND sg13g2_buf_2
XFILLER_103_523 VPWR VGND sg13g2_fill_1
Xplace1696 _07055_ net1696 VPWR VGND sg13g2_buf_2
XFILLER_0_105 VPWR VGND sg13g2_decap_8
Xplace1674 _03453_ net1674 VPWR VGND sg13g2_buf_2
X_09996_ _04083_ VPWR _04084_ VGND _04027_ _04081_ sg13g2_o21ai_1
X_08947_ _03104_ _03133_ _03134_ VPWR VGND sg13g2_nor2_1
XFILLER_103_589 VPWR VGND sg13g2_decap_8
X_08878_ _03023_ _03027_ _03063_ _03064_ _03065_ VPWR VGND sg13g2_nor4_1
XFILLER_57_654 VPWR VGND sg13g2_decap_8
XFILLER_57_632 VPWR VGND sg13g2_decap_8
XFILLER_28_56 VPWR VGND sg13g2_decap_8
X_07829_ _02091_ _02015_ _02125_ VPWR VGND sg13g2_nor2_1
XFILLER_85_985 VPWR VGND sg13g2_decap_8
XFILLER_72_602 VPWR VGND sg13g2_fill_1
XFILLER_57_687 VPWR VGND sg13g2_decap_4
XFILLER_17_518 VPWR VGND sg13g2_decap_4
XFILLER_29_378 VPWR VGND sg13g2_decap_8
XFILLER_84_495 VPWR VGND sg13g2_decap_8
XFILLER_38_890 VPWR VGND sg13g2_decap_8
X_10840_ VPWR _04852_ _04851_ VGND sg13g2_inv_1
XFILLER_72_668 VPWR VGND sg13g2_fill_1
XFILLER_25_551 VPWR VGND sg13g2_decap_8
XFILLER_44_77 VPWR VGND sg13g2_decap_8
X_10771_ fp16_res_pipe.add_renorm0.exp\[7\] net1709 _04783_ VPWR VGND sg13g2_nor2_1
X_13490_ VPWR _00041_ net83 VGND sg13g2_inv_1
X_12510_ fpmul.reg_a_out\[11\] net1953 _06340_ VPWR VGND sg13g2_nor2_1
X_12441_ _06274_ _06273_ _06287_ VPWR VGND sg13g2_and2_1
XFILLER_13_779 VPWR VGND sg13g2_decap_8
XFILLER_40_598 VPWR VGND sg13g2_fill_2
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_21_790 VPWR VGND sg13g2_fill_2
X_12372_ _06195_ _06197_ _06218_ VPWR VGND sg13g2_xor2_1
XFILLER_60_76 VPWR VGND sg13g2_fill_2
XFILLER_125_147 VPWR VGND sg13g2_decap_8
XFILLER_114_0 VPWR VGND sg13g2_decap_8
X_11323_ _03353_ _05026_ _05278_ VPWR VGND sg13g2_nor2_1
X_14111_ VPWR _00662_ net52 VGND sg13g2_inv_1
XFILLER_5_934 VPWR VGND sg13g2_decap_8
Xclkbuf_4_0_0_clk clknet_0_clk clknet_4_0_0_clk VPWR VGND sg13g2_buf_8
XFILLER_109_70 VPWR VGND sg13g2_decap_8
XFILLER_107_851 VPWR VGND sg13g2_decap_8
X_11254_ _05218_ _05217_ net1635 VPWR VGND sg13g2_nand2_1
X_14042_ VPWR _00593_ net20 VGND sg13g2_inv_1
XFILLER_5_49 VPWR VGND sg13g2_decap_8
XFILLER_4_455 VPWR VGND sg13g2_decap_8
XFILLER_106_361 VPWR VGND sg13g2_fill_2
XFILLER_79_223 VPWR VGND sg13g2_decap_8
X_10205_ _04281_ net1830 net1683 fp16_res_pipe.op_sign_logic0.mantisa_b\[8\] _03988_
+ VPWR VGND sg13g2_a22oi_1
XFILLER_122_854 VPWR VGND sg13g2_decap_8
X_11185_ _05154_ net1655 _05073_ VPWR VGND sg13g2_nand2_1
XFILLER_95_738 VPWR VGND sg13g2_decap_8
XFILLER_76_930 VPWR VGND sg13g2_fill_1
X_10136_ _04215_ _04217_ _04218_ VPWR VGND sg13g2_nor2_1
XFILLER_125_91 VPWR VGND sg13g2_decap_8
X_14944_ _00745_ VGND VPWR _01464_ acc_sub.exp_mant_logic0.a\[12\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_1
XFILLER_47_131 VPWR VGND sg13g2_decap_8
X_10067_ _01211_ _04152_ _04154_ VPWR VGND sg13g2_nand2_1
XFILLER_91_922 VPWR VGND sg13g2_decap_8
XFILLER_36_816 VPWR VGND sg13g2_fill_2
XFILLER_91_933 VPWR VGND sg13g2_decap_8
X_14875_ _00676_ VGND VPWR _01395_ acc_sub.exp_mant_logic0.b\[1\] clknet_leaf_58_clk
+ sg13g2_dfrbpq_2
XFILLER_48_698 VPWR VGND sg13g2_fill_2
XFILLER_63_657 VPWR VGND sg13g2_fill_2
XFILLER_51_819 VPWR VGND sg13g2_fill_2
XFILLER_35_359 VPWR VGND sg13g2_decap_8
X_13826_ VPWR _00377_ net10 VGND sg13g2_inv_1
X_13757_ VPWR _00308_ net59 VGND sg13g2_inv_1
XFILLER_44_893 VPWR VGND sg13g2_decap_8
XFILLER_44_882 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_136_clk clknet_5_2__leaf_clk clknet_leaf_136_clk VPWR VGND sg13g2_buf_8
X_10969_ _04969_ _04679_ _04672_ VPWR VGND sg13g2_nand2_1
X_12708_ _06515_ VPWR _00932_ VGND _06510_ _02648_ sg13g2_o21ai_1
XFILLER_43_381 VPWR VGND sg13g2_decap_8
XFILLER_16_595 VPWR VGND sg13g2_fill_2
X_13688_ VPWR _00239_ net59 VGND sg13g2_inv_1
XFILLER_31_576 VPWR VGND sg13g2_fill_2
X_12639_ _06455_ net1851 fpdiv.div_out\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_116_103 VPWR VGND sg13g2_decap_8
X_14309_ _00110_ VGND VPWR _00853_ sipo.bit_counter\[3\] clknet_leaf_6_clk sg13g2_dfrbpq_1
XFILLER_125_681 VPWR VGND sg13g2_decap_8
XFILLER_98_532 VPWR VGND sg13g2_fill_1
XFILLER_113_865 VPWR VGND sg13g2_decap_8
X_09850_ VGND VPWR _03662_ _03840_ _03960_ _03959_ sg13g2_a21oi_1
X_08801_ VPWR _02988_ _02987_ VGND sg13g2_inv_1
X_09781_ _03895_ net1803 _03892_ _03896_ VPWR VGND sg13g2_nand3_1
XFILLER_100_526 VPWR VGND sg13g2_decap_8
XFILLER_100_559 VPWR VGND sg13g2_decap_4
X_08732_ VGND VPWR _01723_ acc_sum.reg1en.d\[0\] _01326_ _02934_ sg13g2_a21oi_1
XFILLER_39_621 VPWR VGND sg13g2_decap_8
XFILLER_22_1003 VPWR VGND sg13g2_decap_8
X_08663_ _02882_ _02738_ _02881_ VPWR VGND sg13g2_xnor2_1
XFILLER_67_985 VPWR VGND sg13g2_decap_8
XFILLER_66_451 VPWR VGND sg13g2_fill_2
XFILLER_39_665 VPWR VGND sg13g2_decap_4
XFILLER_38_142 VPWR VGND sg13g2_fill_1
XFILLER_27_805 VPWR VGND sg13g2_fill_1
XFILLER_82_933 VPWR VGND sg13g2_decap_8
XFILLER_54_646 VPWR VGND sg13g2_decap_4
XFILLER_54_624 VPWR VGND sg13g2_fill_2
XFILLER_53_112 VPWR VGND sg13g2_fill_2
XFILLER_121_49 VPWR VGND sg13g2_decap_8
X_07614_ _01816_ _01909_ _01928_ VPWR VGND sg13g2_nor2_1
X_08594_ _02817_ acc_sum.op_sign_logic0.mantisa_a\[0\] acc_sum.op_sign_logic0.mantisa_b\[0\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_53_156 VPWR VGND sg13g2_decap_8
X_07545_ _01862_ _01779_ acc_sub.seg_reg0.q\[23\] VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_127_clk clknet_5_7__leaf_clk clknet_leaf_127_clk VPWR VGND sg13g2_buf_8
X_07476_ VPWR _01799_ acc_sub.exp_mant_logic0.b\[11\] VGND sg13g2_inv_1
XFILLER_50_841 VPWR VGND sg13g2_decap_8
XFILLER_14_14 VPWR VGND sg13g2_decap_8
XFILLER_22_532 VPWR VGND sg13g2_decap_8
X_09215_ fp16_res_pipe.op_sign_logic0.mantisa_a\[10\] _03368_ _03369_ VPWR VGND sg13g2_nor2_1
X_09146_ net1800 acc_sub.y\[4\] _03322_ VPWR VGND sg13g2_nor2_1
XFILLER_5_219 VPWR VGND sg13g2_decap_4
X_09077_ VGND VPWR net1786 _03260_ _03261_ _03136_ sg13g2_a21oi_1
XFILLER_30_35 VPWR VGND sg13g2_decap_8
XFILLER_123_618 VPWR VGND sg13g2_fill_1
XFILLER_123_607 VPWR VGND sg13g2_decap_8
XFILLER_107_147 VPWR VGND sg13g2_fill_1
X_08028_ _02294_ _02293_ _02185_ VPWR VGND sg13g2_nand2_1
XFILLER_2_926 VPWR VGND sg13g2_decap_8
XFILLER_77_705 VPWR VGND sg13g2_fill_1
XFILLER_1_436 VPWR VGND sg13g2_decap_8
X_09979_ _04068_ VPWR _01213_ VGND _04012_ _04054_ sg13g2_o21ai_1
XFILLER_92_708 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_91_207 VPWR VGND sg13g2_fill_2
XFILLER_58_974 VPWR VGND sg13g2_fill_2
X_12990_ _06758_ _06749_ _06753_ VPWR VGND sg13g2_xnor2_1
XFILLER_57_473 VPWR VGND sg13g2_fill_1
XFILLER_55_21 VPWR VGND sg13g2_decap_8
X_11941_ _05804_ VPWR _00987_ VGND net1874 _05803_ sg13g2_o21ai_1
XFILLER_44_112 VPWR VGND sg13g2_decap_8
XFILLER_29_197 VPWR VGND sg13g2_fill_1
XFILLER_73_966 VPWR VGND sg13g2_decap_8
XFILLER_72_465 VPWR VGND sg13g2_decap_4
XFILLER_55_87 VPWR VGND sg13g2_decap_8
XFILLER_44_156 VPWR VGND sg13g2_fill_1
X_14660_ _00461_ VGND VPWR _01188_ fp16_res_pipe.exp_mant_logic0.b\[13\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
X_11872_ add_result\[2\] _05568_ net1850 _01015_ VPWR VGND sg13g2_mux2_1
XFILLER_72_498 VPWR VGND sg13g2_decap_8
X_13611_ VPWR _00162_ net111 VGND sg13g2_inv_1
XFILLER_60_616 VPWR VGND sg13g2_fill_1
X_14591_ _00392_ VGND VPWR _01123_ fp16_res_pipe.y\[2\] clknet_leaf_128_clk sg13g2_dfrbpq_1
X_10823_ _04835_ _04809_ _04735_ VPWR VGND sg13g2_xnor2_1
Xclkbuf_leaf_118_clk clknet_5_9__leaf_clk clknet_leaf_118_clk VPWR VGND sg13g2_buf_8
X_13542_ VPWR _00093_ net101 VGND sg13g2_inv_1
XFILLER_25_392 VPWR VGND sg13g2_decap_8
XFILLER_71_64 VPWR VGND sg13g2_decap_4
XFILLER_41_863 VPWR VGND sg13g2_decap_8
XFILLER_40_340 VPWR VGND sg13g2_decap_4
X_10754_ _04767_ _04766_ net1822 VPWR VGND sg13g2_nand2_1
X_13473_ VPWR _00024_ net33 VGND sg13g2_inv_1
XFILLER_40_395 VPWR VGND sg13g2_decap_8
XFILLER_9_569 VPWR VGND sg13g2_decap_8
X_10685_ _04698_ _04666_ _04672_ VPWR VGND sg13g2_nand2_1
X_12424_ VPWR _06270_ _06266_ VGND sg13g2_inv_1
XFILLER_127_946 VPWR VGND sg13g2_decap_8
X_12355_ _06201_ _06200_ _06172_ VPWR VGND sg13g2_nand2_1
XFILLER_65_9 VPWR VGND sg13g2_fill_1
XFILLER_5_731 VPWR VGND sg13g2_fill_1
XFILLER_114_618 VPWR VGND sg13g2_decap_4
XFILLER_114_607 VPWR VGND sg13g2_fill_2
XFILLER_99_307 VPWR VGND sg13g2_fill_1
X_11306_ _05264_ net1634 _05263_ VPWR VGND sg13g2_nand2_1
XFILLER_107_681 VPWR VGND sg13g2_fill_1
X_12286_ VPWR _06132_ _06130_ VGND sg13g2_inv_1
X_14025_ VPWR _00576_ net100 VGND sg13g2_inv_1
X_11237_ _05202_ acc_sum.exp_mant_logic0.a\[1\] net1680 acc_sum.op_sign_logic0.mantisa_a\[4\]
+ net1759 VPWR VGND sg13g2_a22oi_1
XFILLER_122_684 VPWR VGND sg13g2_fill_1
XFILLER_121_161 VPWR VGND sg13g2_decap_8
XFILLER_68_716 VPWR VGND sg13g2_decap_8
XFILLER_67_215 VPWR VGND sg13g2_fill_2
XFILLER_110_857 VPWR VGND sg13g2_decap_8
XFILLER_49_952 VPWR VGND sg13g2_fill_2
XFILLER_0_491 VPWR VGND sg13g2_decap_8
X_10119_ _03613_ _04124_ _04202_ VPWR VGND sg13g2_nor2_1
XFILLER_67_259 VPWR VGND sg13g2_decap_8
X_11099_ _02937_ _02939_ _02935_ _05070_ VPWR VGND _02941_ sg13g2_nand4_1
XFILLER_91_730 VPWR VGND sg13g2_decap_8
X_14927_ _00728_ VGND VPWR _01447_ fpdiv.divider0.divisor_reg\[7\] clknet_leaf_85_clk
+ sg13g2_dfrbpq_2
XFILLER_48_473 VPWR VGND sg13g2_decap_8
XFILLER_35_112 VPWR VGND sg13g2_decap_8
XFILLER_91_741 VPWR VGND sg13g2_fill_2
XFILLER_63_465 VPWR VGND sg13g2_decap_8
XFILLER_63_432 VPWR VGND sg13g2_fill_1
X_14858_ _00659_ VGND VPWR _01382_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[9\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_1
X_13809_ VPWR _00360_ net77 VGND sg13g2_inv_1
Xclkbuf_leaf_109_clk clknet_5_10__leaf_clk clknet_leaf_109_clk VPWR VGND sg13g2_buf_8
X_07330_ _01690_ _01692_ _01689_ _01479_ VPWR VGND sg13g2_nand3_1
X_14789_ _00590_ VGND VPWR _01313_ acc_sum.exp_mant_logic0.a\[2\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
XFILLER_50_126 VPWR VGND sg13g2_decap_8
XFILLER_32_841 VPWR VGND sg13g2_decap_8
X_07261_ VGND VPWR _01521_ _01526_ _01631_ _01520_ sg13g2_a21oi_1
X_09000_ acc_sub.add_renorm0.exp\[4\] net1699 _03186_ VPWR VGND sg13g2_nor2_1
XFILLER_31_373 VPWR VGND sg13g2_decap_8
X_07192_ _01561_ _01563_ _01564_ VPWR VGND sg13g2_nor2_2
XFILLER_117_401 VPWR VGND sg13g2_fill_1
XFILLER_77_0 VPWR VGND sg13g2_decap_8
XFILLER_118_957 VPWR VGND sg13g2_decap_8
XFILLER_8_580 VPWR VGND sg13g2_fill_2
XFILLER_117_467 VPWR VGND sg13g2_decap_8
XFILLER_105_618 VPWR VGND sg13g2_fill_1
XFILLER_6_70 VPWR VGND sg13g2_decap_8
XFILLER_104_128 VPWR VGND sg13g2_decap_4
X_09902_ fp16_res_pipe.exp_mant_logic0.b\[13\] _03591_ _03999_ VPWR VGND sg13g2_nor2_1
XFILLER_98_373 VPWR VGND sg13g2_fill_2
X_09833_ _03944_ VPWR _01235_ VGND acc_sum.reg3en.q\[0\] _03934_ sg13g2_o21ai_1
XFILLER_86_524 VPWR VGND sg13g2_decap_8
XFILLER_112_194 VPWR VGND sg13g2_decap_4
XFILLER_86_546 VPWR VGND sg13g2_fill_2
XFILLER_58_237 VPWR VGND sg13g2_fill_1
X_09764_ VGND VPWR _03877_ _03849_ _03880_ _03879_ sg13g2_a21oi_1
X_09695_ _03811_ _02806_ acc_sum.add_renorm0.exp\[3\] VPWR VGND sg13g2_nand2_1
X_08715_ _02924_ acc_sum.add_renorm0.exp\[5\] VPWR VGND sg13g2_inv_2
XFILLER_67_782 VPWR VGND sg13g2_decap_4
XFILLER_27_613 VPWR VGND sg13g2_fill_2
XFILLER_27_635 VPWR VGND sg13g2_fill_1
X_08646_ VPWR _02867_ _02836_ VGND sg13g2_inv_1
XFILLER_70_925 VPWR VGND sg13g2_fill_2
XFILLER_70_914 VPWR VGND sg13g2_decap_8
XFILLER_42_627 VPWR VGND sg13g2_fill_2
XFILLER_25_35 VPWR VGND sg13g2_decap_8
XFILLER_70_958 VPWR VGND sg13g2_decap_8
XFILLER_41_137 VPWR VGND sg13g2_fill_1
XFILLER_41_126 VPWR VGND sg13g2_decap_8
X_07459_ acc_sub.exp_mant_logic0.b\[14\] net1782 _01782_ VPWR VGND sg13g2_nor2_1
XFILLER_50_693 VPWR VGND sg13g2_decap_4
XFILLER_10_524 VPWR VGND sg13g2_decap_8
XFILLER_41_56 VPWR VGND sg13g2_decap_8
X_10470_ _04384_ VPWR _04518_ VGND _04459_ _04456_ sg13g2_o21ai_1
X_09129_ _03160_ _03099_ _03309_ VPWR VGND sg13g2_nor2_1
XFILLER_109_935 VPWR VGND sg13g2_decap_8
X_12140_ VPWR _05986_ _05985_ VGND sg13g2_inv_1
XFILLER_124_949 VPWR VGND sg13g2_decap_8
XFILLER_123_459 VPWR VGND sg13g2_fill_2
XFILLER_89_340 VPWR VGND sg13g2_fill_1
X_12071_ VPWR _05917_ _05916_ VGND sg13g2_inv_1
XFILLER_2_745 VPWR VGND sg13g2_decap_8
XFILLER_1_233 VPWR VGND sg13g2_decap_8
XFILLER_104_673 VPWR VGND sg13g2_decap_8
X_11022_ _04999_ _05000_ _05001_ VPWR VGND sg13g2_nor2_1
XFILLER_49_248 VPWR VGND sg13g2_fill_2
XFILLER_49_237 VPWR VGND sg13g2_fill_1
XFILLER_1_299 VPWR VGND sg13g2_decap_4
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_106_93 VPWR VGND sg13g2_decap_8
XFILLER_66_42 VPWR VGND sg13g2_fill_2
X_12973_ VPWR _06743_ fpmul.reg_p_out\[0\] VGND sg13g2_inv_1
X_14712_ _00513_ VGND VPWR _01240_ acc_sum.y\[15\] clknet_leaf_24_clk sg13g2_dfrbpq_1
X_11924_ VPWR _05793_ fpmul.seg_reg0.q\[38\] VGND sg13g2_inv_1
XFILLER_45_432 VPWR VGND sg13g2_decap_8
XFILLER_122_70 VPWR VGND sg13g2_decap_8
X_14643_ _00444_ VGND VPWR net1835 fp16_res_pipe.reg4en.q\[0\] clknet_leaf_128_clk
+ sg13g2_dfrbpq_1
XFILLER_45_487 VPWR VGND sg13g2_decap_8
XFILLER_18_679 VPWR VGND sg13g2_decap_8
X_11855_ _05753_ net1756 add_result\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_26_690 VPWR VGND sg13g2_decap_8
XFILLER_33_649 VPWR VGND sg13g2_decap_8
XFILLER_41_660 VPWR VGND sg13g2_decap_8
X_11786_ net1757 _05685_ _05688_ _05689_ VPWR VGND sg13g2_nor3_1
XFILLER_14_874 VPWR VGND sg13g2_decap_8
X_14574_ _00375_ VGND VPWR _01106_ fp16_sum_pipe.exp_mant_logic0.b\[1\] clknet_leaf_135_clk
+ sg13g2_dfrbpq_2
X_10806_ VPWR _04818_ _04817_ VGND sg13g2_inv_1
X_13525_ VPWR _00076_ net26 VGND sg13g2_inv_1
XFILLER_9_311 VPWR VGND sg13g2_fill_1
X_10737_ _04716_ _04746_ _04750_ VPWR VGND sg13g2_xor2_1
X_13456_ _07107_ VPWR _00776_ VGND _06929_ net1752 sg13g2_o21ai_1
XFILLER_12_1002 VPWR VGND sg13g2_decap_8
XFILLER_127_743 VPWR VGND sg13g2_decap_8
X_12407_ _06051_ _06024_ _06050_ _06253_ VPWR VGND sg13g2_nand3_1
X_10668_ _04681_ _04621_ _04680_ VPWR VGND sg13g2_xnor2_1
XFILLER_12_1013 VPWR VGND sg13g2_fill_1
XFILLER_126_231 VPWR VGND sg13g2_decap_8
X_13387_ acc_sub.x2\[5\] net1693 _07070_ VPWR VGND sg13g2_nor2_1
X_10599_ _04612_ VPWR _01137_ VGND net1934 _02270_ sg13g2_o21ai_1
XFILLER_115_949 VPWR VGND sg13g2_decap_8
XFILLER_114_404 VPWR VGND sg13g2_fill_1
X_12338_ _06112_ _06111_ _06107_ _06184_ VPWR VGND sg13g2_nand3_1
XFILLER_114_448 VPWR VGND sg13g2_decap_8
X_12269_ VPWR _06115_ _06102_ VGND sg13g2_inv_1
XFILLER_123_960 VPWR VGND sg13g2_decap_8
X_14008_ VPWR _00559_ net19 VGND sg13g2_inv_1
XFILLER_122_470 VPWR VGND sg13g2_decap_8
XFILLER_110_610 VPWR VGND sg13g2_decap_8
XFILLER_96_866 VPWR VGND sg13g2_decap_8
XFILLER_68_557 VPWR VGND sg13g2_decap_8
XFILLER_68_535 VPWR VGND sg13g2_decap_4
XFILLER_96_899 VPWR VGND sg13g2_fill_2
XFILLER_68_568 VPWR VGND sg13g2_decap_8
XFILLER_83_538 VPWR VGND sg13g2_decap_8
XFILLER_49_782 VPWR VGND sg13g2_fill_1
XFILLER_37_966 VPWR VGND sg13g2_decap_8
X_09480_ VGND VPWR _03603_ net1919 _01248_ _03604_ sg13g2_a21oi_1
X_08431_ VPWR _02665_ _02664_ VGND sg13g2_inv_1
XFILLER_63_251 VPWR VGND sg13g2_fill_2
XFILLER_36_487 VPWR VGND sg13g2_decap_8
XFILLER_23_126 VPWR VGND sg13g2_decap_8
X_08362_ _02595_ _02603_ _02605_ VPWR VGND sg13g2_nor2_1
X_07313_ _01677_ net1667 _01627_ VPWR VGND sg13g2_nand2_1
X_08293_ _01364_ _02539_ _02540_ VPWR VGND sg13g2_nand2_1
XFILLER_32_693 VPWR VGND sg13g2_decap_8
X_07244_ _01615_ acc_sub.op_sign_logic0.mantisa_a\[9\] acc_sub.op_sign_logic0.mantisa_b\[9\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_20_899 VPWR VGND sg13g2_decap_8
X_07175_ VPWR _01547_ _01546_ VGND sg13g2_inv_1
XFILLER_118_754 VPWR VGND sg13g2_decap_8
XFILLER_117_231 VPWR VGND sg13g2_decap_8
XFILLER_87_19 VPWR VGND sg13g2_fill_2
XFILLER_120_429 VPWR VGND sg13g2_decap_4
XFILLER_115_1012 VPWR VGND sg13g2_fill_2
XFILLER_114_993 VPWR VGND sg13g2_decap_8
XFILLER_101_621 VPWR VGND sg13g2_decap_8
XFILLER_86_332 VPWR VGND sg13g2_decap_4
XFILLER_59_535 VPWR VGND sg13g2_decap_8
X_09816_ _03817_ _03813_ _03929_ VPWR VGND sg13g2_nor2_1
XFILLER_100_120 VPWR VGND sg13g2_decap_4
XFILLER_87_877 VPWR VGND sg13g2_fill_1
XFILLER_86_343 VPWR VGND sg13g2_decap_8
XFILLER_59_579 VPWR VGND sg13g2_decap_4
X_09747_ _03863_ _03862_ net1690 VPWR VGND sg13g2_nand2_1
XFILLER_86_376 VPWR VGND sg13g2_fill_1
XFILLER_46_218 VPWR VGND sg13g2_decap_8
XFILLER_28_966 VPWR VGND sg13g2_decap_8
X_09678_ net1807 acc_sum.add_renorm0.exp\[7\] _03794_ VPWR VGND sg13g2_nor2_1
XFILLER_70_722 VPWR VGND sg13g2_decap_8
XFILLER_55_796 VPWR VGND sg13g2_decap_8
XFILLER_43_925 VPWR VGND sg13g2_fill_1
XFILLER_43_914 VPWR VGND sg13g2_decap_8
XFILLER_36_56 VPWR VGND sg13g2_decap_8
XFILLER_27_487 VPWR VGND sg13g2_fill_2
X_08629_ VPWR _02851_ _02850_ VGND sg13g2_inv_1
XFILLER_70_788 VPWR VGND sg13g2_fill_2
XFILLER_70_766 VPWR VGND sg13g2_fill_2
XFILLER_35_1013 VPWR VGND sg13g2_fill_1
XFILLER_35_1002 VPWR VGND sg13g2_decap_8
X_11640_ _05545_ _05455_ _05450_ VPWR VGND sg13g2_nand2_1
XFILLER_30_608 VPWR VGND sg13g2_fill_1
XFILLER_11_833 VPWR VGND sg13g2_decap_8
X_11571_ VGND VPWR _05433_ fp16_sum_pipe.add_renorm0.mantisa\[4\] _05476_ fp16_sum_pipe.add_renorm0.mantisa\[5\]
+ sg13g2_a21oi_1
X_13310_ acc\[1\] net1677 _07021_ VPWR VGND sg13g2_nor2_1
X_10522_ _04478_ _04418_ _04563_ VPWR VGND sg13g2_nor2_1
X_14290_ _00091_ VGND VPWR _00834_ acc\[0\] clknet_leaf_50_clk sg13g2_dfrbpq_2
XFILLER_108_253 VPWR VGND sg13g2_decap_4
X_13241_ _06966_ net1729 acc_sum.y\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_6_369 VPWR VGND sg13g2_fill_1
X_10453_ _04501_ _04414_ _04500_ VPWR VGND sg13g2_nand2b_1
XFILLER_10_387 VPWR VGND sg13g2_fill_2
XFILLER_10_398 VPWR VGND sg13g2_fill_2
X_13172_ _06915_ VPWR _00868_ VGND _06914_ _06907_ sg13g2_o21ai_1
X_10384_ _04434_ _04432_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_124_746 VPWR VGND sg13g2_decap_8
XFILLER_123_245 VPWR VGND sg13g2_decap_8
XFILLER_112_908 VPWR VGND sg13g2_decap_8
X_12123_ _05957_ _05960_ _05969_ VPWR VGND sg13g2_nor2_1
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_542 VPWR VGND sg13g2_decap_8
XFILLER_117_70 VPWR VGND sg13g2_decap_8
X_12054_ _05900_ net1856 net1866 VPWR VGND sg13g2_nand2_2
XFILLER_111_429 VPWR VGND sg13g2_decap_8
XFILLER_105_993 VPWR VGND sg13g2_decap_8
XFILLER_104_492 VPWR VGND sg13g2_fill_1
XFILLER_89_170 VPWR VGND sg13g2_fill_1
XFILLER_78_833 VPWR VGND sg13g2_decap_8
XFILLER_77_310 VPWR VGND sg13g2_decap_8
XFILLER_77_52 VPWR VGND sg13g2_decap_4
XFILLER_120_974 VPWR VGND sg13g2_decap_8
XFILLER_93_814 VPWR VGND sg13g2_fill_2
XFILLER_78_866 VPWR VGND sg13g2_decap_8
XFILLER_77_354 VPWR VGND sg13g2_decap_8
XFILLER_77_74 VPWR VGND sg13g2_fill_2
X_11005_ _04988_ VPWR _01107_ VGND net1929 _02468_ sg13g2_o21ai_1
XFILLER_93_847 VPWR VGND sg13g2_decap_8
XFILLER_77_376 VPWR VGND sg13g2_fill_1
XFILLER_65_527 VPWR VGND sg13g2_decap_8
XFILLER_19_922 VPWR VGND sg13g2_decap_8
XFILLER_92_346 VPWR VGND sg13g2_decap_8
XFILLER_58_590 VPWR VGND sg13g2_fill_1
X_12956_ VGND VPWR net1936 add_result\[1\] _06727_ net1950 sg13g2_a21oi_1
XFILLER_19_999 VPWR VGND sg13g2_decap_8
XFILLER_93_95 VPWR VGND sg13g2_decap_4
X_12887_ _06663_ _06662_ net1922 _06664_ VPWR VGND sg13g2_a21o_2
X_11907_ net1880 fpmul.seg_reg0.q\[44\] _05782_ VPWR VGND sg13g2_nor2_1
XFILLER_34_947 VPWR VGND sg13g2_decap_8
XFILLER_33_435 VPWR VGND sg13g2_fill_1
X_14626_ _00427_ VGND VPWR _01158_ fp16_sum_pipe.add_renorm0.exp\[5\] clknet_leaf_98_clk
+ sg13g2_dfrbpq_1
X_11838_ net1837 _05734_ _05732_ _05737_ VPWR VGND _05736_ sg13g2_nand4_1
X_14557_ _00358_ VGND VPWR _01093_ acc_sum.op_sign_logic0.mantisa_a\[9\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
XFILLER_60_298 VPWR VGND sg13g2_fill_2
XFILLER_60_287 VPWR VGND sg13g2_fill_1
XFILLER_42_980 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_40_clk clknet_5_23__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_13508_ VPWR _00059_ net32 VGND sg13g2_inv_1
X_11769_ _05654_ _05672_ _05673_ VPWR VGND sg13g2_nor2_1
X_14488_ _00289_ VGND VPWR _01026_ add_result\[13\] clknet_leaf_99_clk sg13g2_dfrbpq_2
X_13439_ _07098_ VPWR _00784_ VGND _06911_ net1752 sg13g2_o21ai_1
XFILLER_127_562 VPWR VGND sg13g2_decap_8
XFILLER_115_746 VPWR VGND sg13g2_decap_8
XFILLER_6_892 VPWR VGND sg13g2_decap_8
X_08980_ _03166_ _03165_ _03164_ VPWR VGND sg13g2_nand2b_1
XFILLER_114_256 VPWR VGND sg13g2_decap_8
XFILLER_69_822 VPWR VGND sg13g2_decap_8
X_07931_ fp16_sum_pipe.exp_mant_logic0.a\[10\] _02205_ _02206_ VPWR VGND sg13g2_nor2_1
XFILLER_95_140 VPWR VGND sg13g2_decap_8
X_07862_ VPWR _02156_ acc_sub.exp_mant_logic0.b\[1\] VGND sg13g2_inv_1
XFILLER_68_332 VPWR VGND sg13g2_fill_1
XFILLER_113_28 VPWR VGND sg13g2_decap_8
XFILLER_111_985 VPWR VGND sg13g2_decap_8
X_09601_ _03692_ _03697_ _03717_ _03718_ VPWR VGND sg13g2_nor3_1
XFILLER_96_696 VPWR VGND sg13g2_fill_1
XFILLER_69_899 VPWR VGND sg13g2_fill_2
XFILLER_28_207 VPWR VGND sg13g2_decap_8
X_09532_ _03640_ _03630_ _03645_ _03649_ VPWR VGND sg13g2_nor3_2
X_07793_ _02091_ _02048_ _02092_ VPWR VGND sg13g2_nor2_1
XFILLER_37_785 VPWR VGND sg13g2_fill_1
XFILLER_25_903 VPWR VGND sg13g2_decap_8
XFILLER_52_722 VPWR VGND sg13g2_decap_4
XFILLER_51_210 VPWR VGND sg13g2_decap_8
X_09463_ VPWR _03593_ fp16_res_pipe.exp_mant_logic0.a\[12\] VGND sg13g2_inv_1
XFILLER_36_295 VPWR VGND sg13g2_fill_2
XFILLER_36_284 VPWR VGND sg13g2_decap_8
XFILLER_36_273 VPWR VGND sg13g2_fill_1
XFILLER_52_788 VPWR VGND sg13g2_fill_1
XFILLER_52_766 VPWR VGND sg13g2_decap_4
X_09394_ VGND VPWR _03396_ _03539_ _03541_ _03540_ sg13g2_a21oi_1
XFILLER_12_608 VPWR VGND sg13g2_fill_1
X_08345_ _00000_ _00001_ _02588_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_31_clk clknet_5_17__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
XFILLER_20_641 VPWR VGND sg13g2_fill_2
XFILLER_22_14 VPWR VGND sg13g2_decap_8
X_08276_ _02525_ fp16_sum_pipe.exp_mant_logic0.b\[4\] net1658 fp16_sum_pipe.exp_mant_logic0.b\[2\]
+ _02338_ VPWR VGND sg13g2_a22oi_1
X_07227_ _01598_ _01582_ _01597_ VPWR VGND sg13g2_nand2b_1
XFILLER_118_7 VPWR VGND sg13g2_decap_8
X_07158_ VPWR _01530_ _01529_ VGND sg13g2_inv_1
XFILLER_106_702 VPWR VGND sg13g2_fill_2
XFILLER_4_818 VPWR VGND sg13g2_decap_8
XFILLER_3_317 VPWR VGND sg13g2_decap_8
XFILLER_3_339 VPWR VGND sg13g2_fill_1
XFILLER_105_245 VPWR VGND sg13g2_fill_1
XFILLER_79_619 VPWR VGND sg13g2_fill_2
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_121_749 VPWR VGND sg13g2_decap_8
XFILLER_114_790 VPWR VGND sg13g2_decap_8
XFILLER_102_930 VPWR VGND sg13g2_decap_8
XFILLER_99_490 VPWR VGND sg13g2_decap_8
Xfanout131 net140 net131 VPWR VGND sg13g2_buf_2
Xfanout120 net122 net120 VPWR VGND sg13g2_buf_2
XFILLER_59_321 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_98_clk clknet_5_11__leaf_clk clknet_leaf_98_clk VPWR VGND sg13g2_buf_8
XFILLER_120_259 VPWR VGND sg13g2_decap_8
XFILLER_101_440 VPWR VGND sg13g2_decap_8
XFILLER_87_696 VPWR VGND sg13g2_decap_4
XFILLER_47_33 VPWR VGND sg13g2_decap_8
XFILLER_19_207 VPWR VGND sg13g2_fill_2
X_12810_ VPWR _06593_ div_result\[13\] VGND sg13g2_inv_1
XFILLER_28_730 VPWR VGND sg13g2_fill_2
XFILLER_90_839 VPWR VGND sg13g2_decap_8
X_13790_ VPWR _00341_ net20 VGND sg13g2_inv_1
XFILLER_43_711 VPWR VGND sg13g2_decap_8
XFILLER_16_903 VPWR VGND sg13g2_decap_8
XFILLER_27_262 VPWR VGND sg13g2_decap_8
XFILLER_28_763 VPWR VGND sg13g2_fill_2
XFILLER_103_72 VPWR VGND sg13g2_decap_8
X_12741_ _06542_ VPWR _00926_ VGND _06539_ _02648_ sg13g2_o21ai_1
XFILLER_15_424 VPWR VGND sg13g2_decap_8
X_12672_ _06486_ _06416_ _06465_ VPWR VGND sg13g2_xnor2_1
XFILLER_31_928 VPWR VGND sg13g2_decap_8
X_14411_ _00212_ VGND VPWR _00950_ fpmul.reg_a_out\[8\] clknet_leaf_126_clk sg13g2_dfrbpq_2
X_11623_ _05401_ _05415_ _05408_ _05527_ _05528_ VPWR VGND sg13g2_nor4_1
Xclkbuf_leaf_22_clk clknet_5_18__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_8_49 VPWR VGND sg13g2_decap_8
XFILLER_11_641 VPWR VGND sg13g2_fill_2
X_14342_ _00143_ VGND VPWR _00884_ fpmul.reg_p_out\[6\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_10_140 VPWR VGND sg13g2_fill_1
X_11554_ _05458_ _05446_ _05459_ VPWR VGND sg13g2_and2_1
X_11485_ _05395_ VPWR _01034_ VGND net1945 _01763_ sg13g2_o21ai_1
X_14273_ _00074_ VGND VPWR _00824_ fp16_res_pipe.x2\[6\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_6_133 VPWR VGND sg13g2_decap_8
X_10505_ net1848 fp16_sum_pipe.add_renorm0.mantisa\[6\] _04549_ VPWR VGND sg13g2_nor2_1
XFILLER_11_696 VPWR VGND sg13g2_decap_8
XFILLER_7_678 VPWR VGND sg13g2_decap_8
X_10436_ VPWR _04485_ _04484_ VGND sg13g2_inv_1
XFILLER_124_532 VPWR VGND sg13g2_decap_4
XFILLER_3_840 VPWR VGND sg13g2_decap_8
XFILLER_12_91 VPWR VGND sg13g2_decap_8
XFILLER_124_565 VPWR VGND sg13g2_fill_1
XFILLER_98_939 VPWR VGND sg13g2_decap_8
XFILLER_69_107 VPWR VGND sg13g2_decap_8
X_13155_ sipo.bit_counter\[4\] _06900_ _06901_ VPWR VGND sg13g2_nor2_2
X_10367_ VPWR _04417_ _04416_ VGND sg13g2_inv_1
XFILLER_97_427 VPWR VGND sg13g2_fill_1
XFILLER_88_84 VPWR VGND sg13g2_decap_8
X_13086_ _06849_ _06807_ _06763_ VPWR VGND sg13g2_nand2_1
X_12106_ VPWR _05952_ _05890_ VGND sg13g2_inv_1
X_10298_ _04363_ _04365_ _04360_ _04366_ VPWR VGND sg13g2_nand3_1
XFILLER_33_7 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_89_clk clknet_5_24__leaf_clk clknet_leaf_89_clk VPWR VGND sg13g2_buf_8
X_12037_ net1859 net1863 net1858 _05883_ VPWR VGND sg13g2_nand3_1
XFILLER_120_771 VPWR VGND sg13g2_decap_8
XFILLER_78_696 VPWR VGND sg13g2_decap_8
XFILLER_66_836 VPWR VGND sg13g2_decap_8
XFILLER_93_666 VPWR VGND sg13g2_decap_4
XFILLER_93_644 VPWR VGND sg13g2_fill_2
XFILLER_92_121 VPWR VGND sg13g2_fill_2
XFILLER_92_110 VPWR VGND sg13g2_decap_4
XFILLER_66_858 VPWR VGND sg13g2_decap_4
XFILLER_65_346 VPWR VGND sg13g2_decap_8
XFILLER_65_324 VPWR VGND sg13g2_decap_8
X_13988_ VPWR _00539_ net10 VGND sg13g2_inv_1
X_12939_ _06711_ VPWR _06712_ VGND net1962 _06709_ sg13g2_o21ai_1
XFILLER_74_880 VPWR VGND sg13g2_decap_8
XFILLER_46_593 VPWR VGND sg13g2_decap_8
XFILLER_18_273 VPWR VGND sg13g2_fill_2
XFILLER_18_295 VPWR VGND sg13g2_decap_8
XFILLER_61_563 VPWR VGND sg13g2_decap_8
XFILLER_33_232 VPWR VGND sg13g2_fill_1
XFILLER_61_574 VPWR VGND sg13g2_fill_1
XFILLER_15_980 VPWR VGND sg13g2_decap_8
X_14609_ _00410_ VGND VPWR _01141_ fp16_sum_pipe.exp_mant_logic0.a\[4\] clknet_leaf_134_clk
+ sg13g2_dfrbpq_2
XFILLER_105_1000 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_5_6__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_08130_ _01378_ _02390_ _02391_ VPWR VGND sg13g2_nand2_1
XFILLER_21_449 VPWR VGND sg13g2_fill_1
XFILLER_30_983 VPWR VGND sg13g2_decap_8
XFILLER_119_359 VPWR VGND sg13g2_decap_4
X_08061_ _02327_ _02311_ _02326_ VPWR VGND sg13g2_nand2_2
Xplace1801 acc_sub.reg3en.q\[0\] net1801 VPWR VGND sg13g2_buf_2
Xplace1812 acc_sum.exp_mant_logic0.b\[5\] net1812 VPWR VGND sg13g2_buf_2
XFILLER_127_392 VPWR VGND sg13g2_decap_8
XFILLER_115_521 VPWR VGND sg13g2_decap_4
XFILLER_108_28 VPWR VGND sg13g2_decap_8
Xplace1834 net1833 net1834 VPWR VGND sg13g2_buf_1
Xplace1823 fp16_res_pipe.add_renorm0.mantisa\[11\] net1823 VPWR VGND sg13g2_buf_1
Xplace1845 net1844 net1845 VPWR VGND sg13g2_buf_2
Xplace1856 fpmul.reg_a_out\[4\] net1856 VPWR VGND sg13g2_buf_2
Xplace1878 net1877 net1878 VPWR VGND sg13g2_buf_1
Xplace1867 fpmul.reg_b_out\[2\] net1867 VPWR VGND sg13g2_buf_2
X_08963_ VGND VPWR _03148_ _03149_ net1699 _03144_ sg13g2_a21oi_2
XFILLER_102_226 VPWR VGND sg13g2_fill_2
XFILLER_102_215 VPWR VGND sg13g2_decap_8
XFILLER_88_449 VPWR VGND sg13g2_decap_8
Xplace1889 net1885 net1889 VPWR VGND sg13g2_buf_2
XFILLER_25_1001 VPWR VGND sg13g2_decap_8
XFILLER_68_140 VPWR VGND sg13g2_decap_8
XFILLER_25_1012 VPWR VGND sg13g2_fill_2
X_07914_ _02189_ _02186_ fp16_sum_pipe.exp_mant_logic0.b\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_124_49 VPWR VGND sg13g2_decap_8
X_08894_ VGND VPWR _03079_ _03080_ _03081_ net1787 sg13g2_a21oi_1
XFILLER_111_782 VPWR VGND sg13g2_decap_8
XFILLER_96_460 VPWR VGND sg13g2_fill_2
XFILLER_57_814 VPWR VGND sg13g2_decap_8
XFILLER_29_516 VPWR VGND sg13g2_decap_4
X_07845_ _02139_ VPWR _02140_ VGND _02073_ _02015_ sg13g2_o21ai_1
XFILLER_83_110 VPWR VGND sg13g2_decap_8
XFILLER_72_806 VPWR VGND sg13g2_decap_8
XFILLER_56_324 VPWR VGND sg13g2_fill_1
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_29_538 VPWR VGND sg13g2_decap_4
X_07776_ _02077_ net1651 net1795 VPWR VGND sg13g2_nand2_1
XFILLER_84_666 VPWR VGND sg13g2_fill_2
XFILLER_71_349 VPWR VGND sg13g2_decap_8
XFILLER_25_733 VPWR VGND sg13g2_fill_1
X_09446_ _03583_ net1833 fp16_res_pipe.seg_reg0.q\[25\] VPWR VGND sg13g2_nand2_1
XFILLER_12_427 VPWR VGND sg13g2_decap_8
XFILLER_40_747 VPWR VGND sg13g2_fill_2
X_09377_ _03526_ _03382_ _03472_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_35 VPWR VGND sg13g2_decap_8
X_08328_ _02573_ _02571_ _02572_ VPWR VGND sg13g2_nand2_2
X_08259_ _02506_ _02507_ _02508_ _02509_ VPWR VGND sg13g2_nor3_1
XFILLER_20_482 VPWR VGND sg13g2_decap_8
XFILLER_21_994 VPWR VGND sg13g2_decap_8
XFILLER_125_329 VPWR VGND sg13g2_fill_1
XFILLER_4_615 VPWR VGND sg13g2_fill_2
X_11270_ _01086_ _05231_ _05232_ VPWR VGND sg13g2_nand2_1
XFILLER_106_565 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
X_10221_ _04295_ _04294_ net1636 VPWR VGND sg13g2_nand2_1
XFILLER_121_524 VPWR VGND sg13g2_fill_1
XFILLER_106_598 VPWR VGND sg13g2_fill_2
XFILLER_58_21 VPWR VGND sg13g2_fill_1
XFILLER_0_821 VPWR VGND sg13g2_decap_8
X_10152_ _04233_ net1662 _04232_ VPWR VGND sg13g2_nand2_2
X_14960_ _00761_ VGND VPWR _01480_ acc_sub.add_renorm0.mantisa\[4\] clknet_leaf_66_clk
+ sg13g2_dfrbpq_2
X_10083_ _04169_ _04168_ net1637 VPWR VGND sg13g2_nand2_1
XFILLER_75_622 VPWR VGND sg13g2_fill_1
XFILLER_75_611 VPWR VGND sg13g2_decap_8
XFILLER_48_836 VPWR VGND sg13g2_fill_1
X_13911_ VPWR _00462_ net26 VGND sg13g2_inv_1
XFILLER_0_898 VPWR VGND sg13g2_decap_8
X_14891_ _00692_ VGND VPWR _01411_ acc_sub.op_sign_logic0.mantisa_b\[1\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_2
XFILLER_75_633 VPWR VGND sg13g2_decap_8
XFILLER_74_110 VPWR VGND sg13g2_decap_8
XFILLER_75_688 VPWR VGND sg13g2_decap_4
X_13842_ VPWR _00393_ net35 VGND sg13g2_inv_1
XFILLER_90_647 VPWR VGND sg13g2_decap_8
X_13773_ VPWR _00324_ net108 VGND sg13g2_inv_1
XFILLER_28_582 VPWR VGND sg13g2_fill_2
XFILLER_90_669 VPWR VGND sg13g2_fill_2
X_12724_ _06442_ _06528_ _06529_ VPWR VGND sg13g2_nor2_1
X_10985_ _04978_ VPWR _01117_ VGND net1926 _02199_ sg13g2_o21ai_1
XFILLER_15_221 VPWR VGND sg13g2_fill_1
XFILLER_43_574 VPWR VGND sg13g2_decap_8
XFILLER_15_265 VPWR VGND sg13g2_decap_4
X_12655_ _06471_ fpdiv.reg_a_out\[14\] fpdiv.reg_b_out\[14\] VPWR VGND sg13g2_xnor2_1
XFILLER_90_96 VPWR VGND sg13g2_decap_4
X_12586_ _06402_ _06399_ _06401_ VPWR VGND sg13g2_nand2_1
XFILLER_11_460 VPWR VGND sg13g2_fill_2
X_11606_ _05449_ _05444_ _05511_ VPWR VGND sg13g2_nor2_1
X_14325_ _00126_ VGND VPWR _00868_ sipo.word\[13\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_8_965 VPWR VGND sg13g2_decap_8
X_11537_ _05442_ _05440_ _05441_ VPWR VGND sg13g2_nand2_2
XFILLER_125_830 VPWR VGND sg13g2_decap_8
X_11468_ _05386_ VPWR _01042_ VGND net1942 _05385_ sg13g2_o21ai_1
X_14256_ _00057_ VGND VPWR _00807_ acc_sub.x2\[5\] clknet_leaf_17_clk sg13g2_dfrbpq_2
X_11399_ _05344_ net1718 fpdiv.div_out\[6\] VPWR VGND sg13g2_nand2_1
X_14187_ VPWR _00738_ net115 VGND sg13g2_inv_1
X_13207_ VPWR _06939_ sipo.shift_reg\[2\] VGND sg13g2_inv_1
X_10419_ _04459_ _04457_ _04468_ VPWR VGND sg13g2_nor2_1
XFILLER_97_202 VPWR VGND sg13g2_fill_2
X_13138_ _06564_ _06880_ _06556_ _06889_ VPWR VGND sg13g2_nand3_1
XFILLER_3_681 VPWR VGND sg13g2_decap_8
XFILLER_3_692 VPWR VGND sg13g2_fill_1
XFILLER_97_279 VPWR VGND sg13g2_decap_8
XFILLER_78_471 VPWR VGND sg13g2_fill_2
X_13069_ VPWR _06837_ _06835_ VGND sg13g2_inv_1
Xclkbuf_leaf_2_clk clknet_5_1__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_39_847 VPWR VGND sg13g2_decap_8
XFILLER_38_335 VPWR VGND sg13g2_fill_2
X_07630_ VGND VPWR _01932_ _01943_ _01944_ _01855_ sg13g2_a21oi_1
XFILLER_94_975 VPWR VGND sg13g2_decap_8
XFILLER_93_474 VPWR VGND sg13g2_decap_8
XFILLER_66_688 VPWR VGND sg13g2_decap_8
XFILLER_38_379 VPWR VGND sg13g2_fill_1
XFILLER_94_1010 VPWR VGND sg13g2_decap_4
X_07561_ _01874_ VPWR _01875_ VGND _01873_ _01831_ sg13g2_o21ai_1
XFILLER_54_839 VPWR VGND sg13g2_fill_1
XFILLER_0_1003 VPWR VGND sg13g2_decap_8
XFILLER_80_146 VPWR VGND sg13g2_decap_4
X_07492_ acc_sub.exp_mant_logic0.b\[7\] _01739_ _01815_ VPWR VGND sg13g2_nor2_1
XFILLER_34_574 VPWR VGND sg13g2_fill_1
XFILLER_22_725 VPWR VGND sg13g2_decap_8
X_09231_ fp16_res_pipe.op_sign_logic0.mantisa_b\[6\] _03384_ _03385_ VPWR VGND sg13g2_nor2_2
XFILLER_119_112 VPWR VGND sg13g2_decap_8
X_09162_ VPWR _03331_ acc_sum.exp_mant_logic0.b\[13\] VGND sg13g2_inv_1
XFILLER_9_70 VPWR VGND sg13g2_decap_8
X_08113_ _01379_ _02374_ _02375_ VPWR VGND sg13g2_nand2_1
X_09093_ _03196_ _03275_ _03099_ _03276_ VPWR VGND sg13g2_a21o_1
XFILLER_119_49 VPWR VGND sg13g2_decap_8
XFILLER_119_189 VPWR VGND sg13g2_decap_8
X_08044_ VGND VPWR _02231_ _02245_ _02310_ _02309_ sg13g2_a21oi_1
XFILLER_116_863 VPWR VGND sg13g2_decap_8
Xplace1653 _05181_ net1653 VPWR VGND sg13g2_buf_2
Xplace1642 _04190_ net1642 VPWR VGND sg13g2_buf_1
Xplace1664 _03681_ net1664 VPWR VGND sg13g2_buf_2
XFILLER_103_535 VPWR VGND sg13g2_fill_1
Xplace1686 _01840_ net1686 VPWR VGND sg13g2_buf_2
XFILLER_89_725 VPWR VGND sg13g2_decap_8
Xplace1675 _03453_ net1675 VPWR VGND sg13g2_buf_2
Xplace1697 _05075_ net1697 VPWR VGND sg13g2_buf_1
X_09995_ VGND VPWR _04082_ _04019_ _04083_ _04033_ sg13g2_a21oi_1
X_08946_ _03120_ _03125_ _03113_ _03133_ VPWR VGND _03132_ sg13g2_nand4_1
XFILLER_88_279 VPWR VGND sg13g2_decap_8
XFILLER_57_600 VPWR VGND sg13g2_decap_8
X_08877_ _03064_ _03034_ _03038_ VPWR VGND sg13g2_nand2_1
XFILLER_85_964 VPWR VGND sg13g2_decap_8
XFILLER_28_35 VPWR VGND sg13g2_decap_8
XFILLER_29_335 VPWR VGND sg13g2_fill_2
X_07828_ _02073_ _01977_ _02124_ VPWR VGND sg13g2_nor2_1
XFILLER_71_113 VPWR VGND sg13g2_decap_8
X_07759_ VPWR _02062_ _01847_ VGND sg13g2_inv_1
XFILLER_71_146 VPWR VGND sg13g2_fill_1
XFILLER_25_530 VPWR VGND sg13g2_decap_8
XFILLER_25_541 VPWR VGND sg13g2_fill_1
XFILLER_44_56 VPWR VGND sg13g2_decap_8
XFILLER_40_500 VPWR VGND sg13g2_decap_8
X_10770_ _04782_ _03574_ _04781_ VPWR VGND sg13g2_xnor2_1
XFILLER_13_725 VPWR VGND sg13g2_fill_2
X_09429_ _03571_ VPWR _01266_ VGND fp16_res_pipe.reg2en.q\[0\] _03565_ sg13g2_o21ai_1
XFILLER_9_707 VPWR VGND sg13g2_fill_1
XFILLER_13_758 VPWR VGND sg13g2_fill_2
XFILLER_25_596 VPWR VGND sg13g2_fill_2
X_12440_ VGND VPWR _06267_ _06272_ _06286_ _06285_ sg13g2_a21oi_1
XFILLER_40_577 VPWR VGND sg13g2_decap_8
XFILLER_21_780 VPWR VGND sg13g2_decap_8
X_12371_ _06217_ _06213_ _06216_ VPWR VGND sg13g2_nand2_1
XFILLER_60_88 VPWR VGND sg13g2_decap_8
X_14110_ VPWR _00661_ net52 VGND sg13g2_inv_1
XFILLER_5_913 VPWR VGND sg13g2_decap_8
XFILLER_125_126 VPWR VGND sg13g2_decap_8
X_11322_ _03347_ _05143_ _05277_ VPWR VGND sg13g2_nor2_1
XFILLER_60_99 VPWR VGND sg13g2_fill_1
XFILLER_5_28 VPWR VGND sg13g2_decap_8
XFILLER_4_434 VPWR VGND sg13g2_decap_8
XFILLER_107_0 VPWR VGND sg13g2_decap_4
XFILLER_106_340 VPWR VGND sg13g2_decap_8
X_14041_ VPWR _00592_ net76 VGND sg13g2_inv_1
X_11253_ _05208_ _05216_ _05207_ _05217_ VPWR VGND sg13g2_nand3_1
XFILLER_122_833 VPWR VGND sg13g2_decap_8
XFILLER_69_53 VPWR VGND sg13g2_fill_1
X_10204_ _04280_ net1636 _04279_ VPWR VGND sg13g2_nand2_1
XFILLER_121_343 VPWR VGND sg13g2_decap_4
XFILLER_125_70 VPWR VGND sg13g2_decap_8
XFILLER_79_279 VPWR VGND sg13g2_fill_2
XFILLER_76_920 VPWR VGND sg13g2_decap_4
XFILLER_48_611 VPWR VGND sg13g2_fill_1
XFILLER_0_651 VPWR VGND sg13g2_decap_8
X_10135_ _04216_ VPWR _04217_ VGND _03617_ net1703 sg13g2_o21ai_1
XFILLER_102_590 VPWR VGND sg13g2_decap_8
X_14943_ _00744_ VGND VPWR _01463_ acc_sub.exp_mant_logic0.a\[11\] clknet_leaf_51_clk
+ sg13g2_dfrbpq_1
XFILLER_47_110 VPWR VGND sg13g2_decap_8
XFILLER_0_684 VPWR VGND sg13g2_decap_8
X_10066_ _04154_ net1827 net1682 fp16_res_pipe.op_sign_logic0.mantisa_a\[9\] net1764
+ VPWR VGND sg13g2_a22oi_1
X_14874_ _00675_ VGND VPWR _01394_ acc_sub.exp_mant_logic0.b\[0\] clknet_leaf_59_clk
+ sg13g2_dfrbpq_2
XFILLER_85_85 VPWR VGND sg13g2_decap_8
XFILLER_75_463 VPWR VGND sg13g2_decap_8
XFILLER_90_400 VPWR VGND sg13g2_fill_1
XFILLER_85_96 VPWR VGND sg13g2_decap_8
XFILLER_75_496 VPWR VGND sg13g2_fill_1
XFILLER_75_474 VPWR VGND sg13g2_fill_1
XFILLER_35_338 VPWR VGND sg13g2_fill_2
X_13825_ VPWR _00376_ net10 VGND sg13g2_inv_1
XFILLER_91_989 VPWR VGND sg13g2_decap_8
XFILLER_44_861 VPWR VGND sg13g2_decap_8
X_13756_ VPWR _00307_ net108 VGND sg13g2_inv_1
X_10968_ _04968_ _04670_ _04695_ VPWR VGND sg13g2_nand2_1
XFILLER_16_574 VPWR VGND sg13g2_fill_2
XFILLER_31_511 VPWR VGND sg13g2_decap_4
X_12707_ _06513_ VPWR _06515_ VGND net1734 _06512_ sg13g2_o21ai_1
X_13687_ VPWR _00238_ net61 VGND sg13g2_inv_1
X_12638_ _06454_ _06421_ _05337_ VPWR VGND sg13g2_nand2_1
X_10899_ VGND VPWR _04889_ _04908_ _04909_ _04742_ sg13g2_a21oi_1
X_12569_ _06385_ fpdiv.reg_a_out\[10\] fpdiv.reg_b_out\[10\] VPWR VGND sg13g2_xnor2_1
X_14308_ _00109_ VGND VPWR _00852_ sipo.bit_counter\[2\] clknet_leaf_8_clk sg13g2_dfrbpq_1
XFILLER_7_261 VPWR VGND sg13g2_decap_4
XFILLER_116_159 VPWR VGND sg13g2_decap_8
X_14239_ _00040_ VGND VPWR _00790_ instr\[4\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_98_500 VPWR VGND sg13g2_decap_8
X_08800_ _02969_ _02986_ _02987_ VPWR VGND sg13g2_nor2_1
XFILLER_113_844 VPWR VGND sg13g2_decap_8
XFILLER_86_706 VPWR VGND sg13g2_decap_8
XFILLER_112_365 VPWR VGND sg13g2_decap_8
X_09780_ _03895_ _03663_ _03894_ _03893_ _03648_ VPWR VGND sg13g2_a22oi_1
XFILLER_85_205 VPWR VGND sg13g2_fill_2
XFILLER_22_0 VPWR VGND sg13g2_decap_8
X_08731_ acc_sum.exp_mant_logic0.a\[15\] acc_sum.reg1en.d\[0\] _02934_ VPWR VGND sg13g2_nor2_1
XFILLER_66_430 VPWR VGND sg13g2_decap_8
X_08662_ _02832_ VPWR _02881_ VGND net1740 _02880_ sg13g2_o21ai_1
XFILLER_82_912 VPWR VGND sg13g2_decap_8
XFILLER_67_975 VPWR VGND sg13g2_decap_4
X_07613_ _01818_ _01913_ _01919_ _01927_ VPWR VGND sg13g2_nand3_1
XFILLER_27_839 VPWR VGND sg13g2_decap_8
XFILLER_121_28 VPWR VGND sg13g2_decap_8
XFILLER_82_989 VPWR VGND sg13g2_decap_8
XFILLER_81_433 VPWR VGND sg13g2_decap_8
X_08593_ _02816_ _02760_ _02764_ VPWR VGND sg13g2_nand2_2
XFILLER_54_658 VPWR VGND sg13g2_decap_4
X_07544_ _01861_ _01847_ acc_sub.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_81_499 VPWR VGND sg13g2_decap_4
XFILLER_22_500 VPWR VGND sg13g2_decap_8
X_07475_ acc_sub.exp_mant_logic0.b\[11\] _01731_ _01798_ VPWR VGND sg13g2_nor2_1
X_09214_ VPWR _03368_ fp16_res_pipe.op_sign_logic0.mantisa_b\[10\] VGND sg13g2_inv_1
XFILLER_22_555 VPWR VGND sg13g2_decap_8
XFILLER_22_566 VPWR VGND sg13g2_fill_2
XFILLER_22_599 VPWR VGND sg13g2_decap_8
XFILLER_108_627 VPWR VGND sg13g2_fill_1
X_09145_ VGND VPWR _03046_ net1801 _01300_ _03321_ sg13g2_a21oi_1
XFILLER_30_14 VPWR VGND sg13g2_decap_8
X_09076_ _03260_ _03236_ _03234_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_905 VPWR VGND sg13g2_decap_8
X_08027_ _02292_ VPWR _02293_ VGND _02245_ _02287_ sg13g2_o21ai_1
XFILLER_116_693 VPWR VGND sg13g2_decap_8
XFILLER_104_833 VPWR VGND sg13g2_decap_8
XFILLER_89_511 VPWR VGND sg13g2_decap_8
XFILLER_1_415 VPWR VGND sg13g2_decap_8
XFILLER_103_321 VPWR VGND sg13g2_fill_1
XFILLER_39_56 VPWR VGND sg13g2_decap_8
X_09978_ _04068_ fp16_res_pipe.exp_mant_logic0.a\[7\] _04056_ net1765 fp16_res_pipe.seg_reg0.q\[22\]
+ VPWR VGND sg13g2_a22oi_1
X_08929_ _03116_ _03017_ _03001_ VPWR VGND sg13g2_nand2_1
XFILLER_73_901 VPWR VGND sg13g2_fill_1
XFILLER_58_964 VPWR VGND sg13g2_fill_2
X_11940_ _05804_ net1877 fpmul.reg_b_out\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_72_411 VPWR VGND sg13g2_fill_2
XFILLER_57_485 VPWR VGND sg13g2_decap_4
XFILLER_45_636 VPWR VGND sg13g2_fill_1
XFILLER_45_614 VPWR VGND sg13g2_decap_8
XFILLER_18_828 VPWR VGND sg13g2_decap_8
XFILLER_72_444 VPWR VGND sg13g2_decap_8
X_11871_ VGND VPWR _05562_ net1850 _01016_ _05763_ sg13g2_a21oi_1
XFILLER_26_850 VPWR VGND sg13g2_fill_1
X_13610_ VPWR _00161_ net111 VGND sg13g2_inv_1
X_14590_ _00391_ VGND VPWR _01122_ fp16_res_pipe.y\[1\] clknet_leaf_127_clk sg13g2_dfrbpq_1
XFILLER_32_319 VPWR VGND sg13g2_decap_8
X_10822_ net1772 _04821_ _04833_ _04834_ VPWR VGND sg13g2_nor3_1
X_13541_ VPWR _00092_ net90 VGND sg13g2_inv_1
X_10753_ _04764_ _04765_ _04763_ _04766_ VPWR VGND sg13g2_nand3_1
XFILLER_25_371 VPWR VGND sg13g2_fill_2
XFILLER_71_43 VPWR VGND sg13g2_decap_4
XFILLER_9_526 VPWR VGND sg13g2_decap_4
X_13472_ VPWR _00023_ net82 VGND sg13g2_inv_1
X_10684_ _04697_ _04675_ _04679_ net1710 _04647_ VPWR VGND sg13g2_a22oi_1
XFILLER_127_925 VPWR VGND sg13g2_decap_8
XFILLER_126_402 VPWR VGND sg13g2_decap_4
X_12423_ _06269_ net1864 _06255_ VPWR VGND sg13g2_nand2b_1
X_12354_ _06200_ _06199_ _06158_ VPWR VGND sg13g2_nand2b_1
XFILLER_126_457 VPWR VGND sg13g2_decap_4
X_11305_ _05261_ _05262_ _05260_ _05263_ VPWR VGND sg13g2_nand3_1
XFILLER_4_231 VPWR VGND sg13g2_fill_2
X_14024_ VPWR _00575_ net98 VGND sg13g2_inv_1
X_12285_ _06131_ _06127_ _06130_ VPWR VGND sg13g2_nand2_1
XFILLER_4_264 VPWR VGND sg13g2_decap_4
X_11236_ _05201_ _05200_ net1635 VPWR VGND sg13g2_nand2_1
XFILLER_45_1004 VPWR VGND sg13g2_decap_8
XFILLER_121_140 VPWR VGND sg13g2_decap_8
XFILLER_95_514 VPWR VGND sg13g2_fill_1
X_11167_ net1663 _05135_ _05136_ VPWR VGND sg13g2_nor2b_1
XFILLER_110_836 VPWR VGND sg13g2_decap_8
XFILLER_96_84 VPWR VGND sg13g2_decap_4
XFILLER_67_227 VPWR VGND sg13g2_decap_8
XFILLER_49_931 VPWR VGND sg13g2_decap_8
XFILLER_0_470 VPWR VGND sg13g2_decap_8
X_10118_ _03605_ _04189_ _04201_ VPWR VGND sg13g2_nor2_1
X_11098_ _02945_ _02947_ _02943_ _05069_ VPWR VGND _02949_ sg13g2_nand4_1
XFILLER_48_452 VPWR VGND sg13g2_decap_8
X_14926_ _00727_ VGND VPWR _01446_ fpdiv.divider0.divisor_reg\[6\] clknet_leaf_75_clk
+ sg13g2_dfrbpq_1
XFILLER_64_934 VPWR VGND sg13g2_decap_4
XFILLER_48_485 VPWR VGND sg13g2_decap_8
X_10049_ VPWR _04137_ _04016_ VGND sg13g2_inv_1
XFILLER_35_135 VPWR VGND sg13g2_decap_8
X_14857_ _00658_ VGND VPWR _01381_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[8\] clknet_5_8__leaf_clk
+ sg13g2_dfrbpq_1
X_13808_ VPWR _00359_ net81 VGND sg13g2_inv_1
X_14788_ _00589_ VGND VPWR _01312_ acc_sum.exp_mant_logic0.a\[1\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_2
XFILLER_64_989 VPWR VGND sg13g2_decap_8
XFILLER_63_488 VPWR VGND sg13g2_decap_8
XFILLER_51_628 VPWR VGND sg13g2_decap_8
XFILLER_50_105 VPWR VGND sg13g2_decap_8
XFILLER_90_285 VPWR VGND sg13g2_fill_2
X_13739_ VPWR _00290_ net55 VGND sg13g2_inv_1
XFILLER_52_1008 VPWR VGND sg13g2_decap_4
XFILLER_31_352 VPWR VGND sg13g2_decap_8
X_07260_ VPWR _01630_ _01629_ VGND sg13g2_inv_1
XFILLER_31_396 VPWR VGND sg13g2_decap_4
X_07191_ acc_sub.op_sign_logic0.mantisa_b\[2\] _01562_ _01563_ VPWR VGND sg13g2_nor2_1
XFILLER_118_936 VPWR VGND sg13g2_decap_8
XFILLER_117_446 VPWR VGND sg13g2_decap_8
X_09901_ VPWR _03998_ _03997_ VGND sg13g2_inv_1
XFILLER_113_674 VPWR VGND sg13g2_decap_8
XFILLER_101_825 VPWR VGND sg13g2_decap_8
X_09832_ _03783_ _03943_ _03941_ _03944_ VPWR VGND sg13g2_nand3_1
X_09763_ _03840_ _03878_ _03879_ VPWR VGND sg13g2_nor2_1
XFILLER_112_162 VPWR VGND sg13g2_decap_8
XFILLER_101_836 VPWR VGND sg13g2_fill_1
XFILLER_100_335 VPWR VGND sg13g2_decap_4
X_08714_ VGND VPWR net1814 _02922_ _01333_ _02923_ sg13g2_a21oi_1
XFILLER_86_569 VPWR VGND sg13g2_decap_8
XFILLER_67_761 VPWR VGND sg13g2_decap_8
XFILLER_39_441 VPWR VGND sg13g2_fill_2
X_09694_ _03810_ _02926_ _03788_ VPWR VGND sg13g2_xnor2_1
XFILLER_73_219 VPWR VGND sg13g2_decap_8
XFILLER_55_923 VPWR VGND sg13g2_decap_4
XFILLER_26_102 VPWR VGND sg13g2_fill_2
X_08645_ _02724_ VPWR _02866_ VGND _02864_ _02865_ sg13g2_o21ai_1
XFILLER_70_904 VPWR VGND sg13g2_decap_4
XFILLER_55_956 VPWR VGND sg13g2_decap_4
XFILLER_15_809 VPWR VGND sg13g2_fill_1
XFILLER_27_658 VPWR VGND sg13g2_decap_4
X_08576_ VGND VPWR _02798_ _02800_ _02799_ _02794_ sg13g2_a21oi_2
XFILLER_81_252 VPWR VGND sg13g2_decap_8
XFILLER_42_606 VPWR VGND sg13g2_decap_8
XFILLER_41_105 VPWR VGND sg13g2_decap_8
XFILLER_25_14 VPWR VGND sg13g2_decap_8
XFILLER_42_639 VPWR VGND sg13g2_decap_4
XFILLER_34_190 VPWR VGND sg13g2_decap_4
XFILLER_23_864 VPWR VGND sg13g2_fill_1
XFILLER_109_914 VPWR VGND sg13g2_decap_8
X_07389_ _01734_ VPWR _01462_ VGND net1893 _01733_ sg13g2_o21ai_1
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_10_569 VPWR VGND sg13g2_fill_2
X_09128_ _03161_ _03096_ _03308_ VPWR VGND sg13g2_nor2_1
XFILLER_124_928 VPWR VGND sg13g2_decap_8
XFILLER_123_427 VPWR VGND sg13g2_decap_8
XFILLER_117_991 VPWR VGND sg13g2_decap_8
X_09059_ _03244_ acc_sub.y\[13\] VPWR VGND sg13g2_inv_2
XFILLER_2_724 VPWR VGND sg13g2_decap_8
XFILLER_89_330 VPWR VGND sg13g2_fill_1
X_12070_ _05916_ net1856 net1864 VPWR VGND sg13g2_nand2_1
XFILLER_104_652 VPWR VGND sg13g2_decap_8
XFILLER_103_140 VPWR VGND sg13g2_fill_2
X_11021_ acc_sum.exp_mant_logic0.a\[12\] _03333_ _05000_ VPWR VGND sg13g2_nor2_2
XFILLER_1_256 VPWR VGND sg13g2_fill_2
XFILLER_106_50 VPWR VGND sg13g2_decap_4
XFILLER_77_525 VPWR VGND sg13g2_decap_8
XFILLER_49_227 VPWR VGND sg13g2_fill_1
XFILLER_92_506 VPWR VGND sg13g2_fill_2
XFILLER_77_558 VPWR VGND sg13g2_decap_4
XFILLER_66_21 VPWR VGND sg13g2_decap_8
XFILLER_65_709 VPWR VGND sg13g2_fill_2
XFILLER_100_891 VPWR VGND sg13g2_fill_2
XFILLER_92_517 VPWR VGND sg13g2_fill_1
X_12972_ _06742_ _06738_ _06741_ _06539_ net1949 VPWR VGND sg13g2_a22oi_1
X_14711_ _00512_ VGND VPWR _01239_ acc_sum.y\[14\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_72_230 VPWR VGND sg13g2_fill_1
XFILLER_46_978 VPWR VGND sg13g2_fill_1
X_11923_ _05792_ VPWR _00993_ VGND net1882 _05791_ sg13g2_o21ai_1
XFILLER_18_658 VPWR VGND sg13g2_decap_8
XFILLER_73_786 VPWR VGND sg13g2_decap_8
XFILLER_72_263 VPWR VGND sg13g2_decap_8
X_14642_ _00443_ VGND VPWR _01174_ fp16_sum_pipe.seg_reg1.q\[21\] clknet_leaf_111_clk
+ sg13g2_dfrbpq_2
X_11854_ _05748_ _05751_ _05570_ _05752_ VPWR VGND sg13g2_nand3_1
XFILLER_33_628 VPWR VGND sg13g2_decap_8
XFILLER_82_53 VPWR VGND sg13g2_fill_1
XFILLER_82_42 VPWR VGND sg13g2_decap_8
XFILLER_72_274 VPWR VGND sg13g2_fill_1
XFILLER_45_499 VPWR VGND sg13g2_decap_8
X_10805_ VGND VPWR _04816_ _04817_ _04815_ net1709 sg13g2_a21oi_2
XFILLER_32_127 VPWR VGND sg13g2_fill_1
X_11785_ VGND VPWR _05687_ _05629_ _05688_ _05495_ sg13g2_a21oi_1
X_14573_ _00374_ VGND VPWR _01105_ fp16_sum_pipe.exp_mant_logic0.b\[0\] clknet_leaf_116_clk
+ sg13g2_dfrbpq_2
XFILLER_14_853 VPWR VGND sg13g2_decap_8
X_13524_ VPWR _00075_ net84 VGND sg13g2_inv_1
XFILLER_9_323 VPWR VGND sg13g2_decap_4
XFILLER_13_363 VPWR VGND sg13g2_decap_4
X_10736_ _04746_ _04630_ _04749_ VPWR VGND sg13g2_nor2_1
X_13455_ _07107_ net1752 sipo.shift_reg\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_40_182 VPWR VGND sg13g2_decap_8
X_10667_ _04641_ fp16_res_pipe.add_renorm0.mantisa\[4\] _04680_ VPWR VGND sg13g2_nor2b_1
XFILLER_127_722 VPWR VGND sg13g2_decap_8
XFILLER_126_210 VPWR VGND sg13g2_decap_8
X_12406_ _06252_ _06148_ _06251_ VPWR VGND sg13g2_nand2_1
X_13386_ _07069_ VPWR _00808_ VGND _06346_ net1694 sg13g2_o21ai_1
X_10598_ _04612_ acc_sub.x2\[0\] net1933 VPWR VGND sg13g2_nand2_1
XFILLER_127_799 VPWR VGND sg13g2_decap_8
XFILLER_126_287 VPWR VGND sg13g2_decap_8
XFILLER_115_928 VPWR VGND sg13g2_decap_8
X_12337_ _06183_ _06182_ _06110_ VPWR VGND sg13g2_nand2_1
XFILLER_5_551 VPWR VGND sg13g2_decap_8
XFILLER_114_438 VPWR VGND sg13g2_fill_1
X_12268_ VGND VPWR _06107_ _06111_ _06114_ _06113_ sg13g2_a21oi_1
XFILLER_68_514 VPWR VGND sg13g2_decap_8
X_11219_ _02953_ _05143_ _05185_ VPWR VGND sg13g2_nor2_1
X_14007_ VPWR _00558_ net19 VGND sg13g2_inv_1
XFILLER_96_845 VPWR VGND sg13g2_decap_8
X_12199_ VGND VPWR _06001_ _05987_ _06045_ _06044_ sg13g2_a21oi_1
XFILLER_64_720 VPWR VGND sg13g2_decap_8
XFILLER_48_271 VPWR VGND sg13g2_fill_1
X_14909_ _00710_ VGND VPWR _01429_ acc_sub.op_sign_logic0.mantisa_a\[8\] clknet_leaf_62_clk
+ sg13g2_dfrbpq_1
XFILLER_63_230 VPWR VGND sg13g2_decap_8
XFILLER_37_945 VPWR VGND sg13g2_decap_8
XFILLER_36_422 VPWR VGND sg13g2_decap_8
X_08430_ _02664_ _02661_ _02663_ VPWR VGND sg13g2_nand2_1
XFILLER_91_572 VPWR VGND sg13g2_decap_8
XFILLER_63_296 VPWR VGND sg13g2_fill_1
XFILLER_51_447 VPWR VGND sg13g2_decap_8
XFILLER_16_190 VPWR VGND sg13g2_decap_8
X_07312_ _01676_ VPWR _01481_ VGND _01656_ _01674_ sg13g2_o21ai_1
XFILLER_60_981 VPWR VGND sg13g2_decap_8
X_08292_ _02540_ net1778 fp16_sum_pipe.op_sign_logic0.mantisa_b\[2\] VPWR VGND sg13g2_nand2_1
X_07243_ _01614_ _01613_ _01514_ VPWR VGND sg13g2_nand2_1
XFILLER_20_856 VPWR VGND sg13g2_decap_8
XFILLER_20_867 VPWR VGND sg13g2_fill_1
XFILLER_31_193 VPWR VGND sg13g2_decap_4
XFILLER_118_733 VPWR VGND sg13g2_decap_8
XFILLER_117_210 VPWR VGND sg13g2_decap_8
X_07174_ acc_sub.op_sign_logic0.mantisa_a\[0\] _01545_ _01546_ VPWR VGND sg13g2_nor2_1
XFILLER_11_49 VPWR VGND sg13g2_decap_8
XFILLER_127_49 VPWR VGND sg13g2_decap_8
XFILLER_120_419 VPWR VGND sg13g2_fill_2
XFILLER_114_972 VPWR VGND sg13g2_decap_8
XFILLER_99_672 VPWR VGND sg13g2_decap_4
XFILLER_99_661 VPWR VGND sg13g2_fill_2
X_09815_ _03927_ net1803 _03928_ VPWR VGND _03924_ sg13g2_nand3b_1
XFILLER_87_823 VPWR VGND sg13g2_decap_8
XFILLER_86_311 VPWR VGND sg13g2_decap_8
XFILLER_59_525 VPWR VGND sg13g2_fill_2
XFILLER_87_867 VPWR VGND sg13g2_decap_8
XFILLER_59_558 VPWR VGND sg13g2_decap_8
XFILLER_101_699 VPWR VGND sg13g2_fill_1
X_09746_ VPWR _03862_ _03793_ VGND sg13g2_inv_1
X_09677_ _03793_ _02920_ _03792_ VPWR VGND sg13g2_xnor2_1
XFILLER_67_591 VPWR VGND sg13g2_fill_1
XFILLER_55_742 VPWR VGND sg13g2_decap_8
XFILLER_36_35 VPWR VGND sg13g2_decap_8
XFILLER_27_422 VPWR VGND sg13g2_decap_8
XFILLER_28_945 VPWR VGND sg13g2_decap_8
X_08628_ VGND VPWR _02849_ _02774_ _02850_ _02773_ sg13g2_a21oi_1
XFILLER_55_775 VPWR VGND sg13g2_decap_8
XFILLER_54_274 VPWR VGND sg13g2_decap_4
XFILLER_43_959 VPWR VGND sg13g2_decap_8
XFILLER_27_499 VPWR VGND sg13g2_decap_4
X_08559_ VPWR _02783_ _02771_ VGND sg13g2_inv_1
XFILLER_11_812 VPWR VGND sg13g2_fill_1
X_11570_ _05475_ _05474_ VPWR VGND sg13g2_inv_2
XFILLER_52_67 VPWR VGND sg13g2_fill_1
X_10521_ VPWR _04562_ _04481_ VGND sg13g2_inv_1
X_13240_ _06965_ net1711 acc_sub.y\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_11_889 VPWR VGND sg13g2_decap_8
XFILLER_109_755 VPWR VGND sg13g2_decap_8
X_10452_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[0\] _04413_ _04500_ VPWR VGND sg13g2_nor2_1
XFILLER_124_725 VPWR VGND sg13g2_decap_8
XFILLER_124_703 VPWR VGND sg13g2_decap_8
X_13171_ _06915_ _06907_ sipo.word\[13\] VPWR VGND sg13g2_nand2_1
X_10383_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[4\] _04432_ _04433_ VPWR VGND sg13g2_nor2_2
XFILLER_123_224 VPWR VGND sg13g2_decap_8
XFILLER_108_298 VPWR VGND sg13g2_decap_8
X_12122_ _05902_ _05967_ _05968_ VPWR VGND sg13g2_nor2_1
XFILLER_2_521 VPWR VGND sg13g2_decap_8
XFILLER_111_408 VPWR VGND sg13g2_fill_1
XFILLER_105_972 VPWR VGND sg13g2_decap_8
X_12053_ _05899_ net1855 net1865 VPWR VGND sg13g2_nand2_2
X_11004_ _04988_ fp16_res_pipe.x2\[2\] net1927 VPWR VGND sg13g2_nand2_1
XFILLER_120_953 VPWR VGND sg13g2_decap_8
XFILLER_78_889 VPWR VGND sg13g2_fill_1
XFILLER_77_86 VPWR VGND sg13g2_fill_1
XFILLER_19_901 VPWR VGND sg13g2_decap_8
X_12955_ _00007_ net1731 net1702 _06726_ VPWR VGND sg13g2_nand3_1
XFILLER_46_720 VPWR VGND sg13g2_decap_4
XFILLER_18_422 VPWR VGND sg13g2_fill_2
XFILLER_93_52 VPWR VGND sg13g2_fill_2
X_11906_ _05781_ fpmul.reg_a_out\[5\] VPWR VGND sg13g2_inv_2
XFILLER_34_926 VPWR VGND sg13g2_decap_8
XFILLER_18_477 VPWR VGND sg13g2_decap_8
XFILLER_19_978 VPWR VGND sg13g2_decap_8
XFILLER_73_594 VPWR VGND sg13g2_decap_8
X_12886_ _06663_ net1909 fp16_res_pipe.y\[7\] VPWR VGND sg13g2_nand2_1
X_14625_ _00426_ VGND VPWR _01157_ fp16_sum_pipe.add_renorm0.exp\[4\] clknet_leaf_120_clk
+ sg13g2_dfrbpq_1
XFILLER_14_650 VPWR VGND sg13g2_fill_2
XFILLER_21_609 VPWR VGND sg13g2_fill_2
X_11837_ _05496_ _05735_ _05736_ VPWR VGND _05619_ sg13g2_nand3b_1
X_14556_ _00357_ VGND VPWR _01092_ acc_sum.op_sign_logic0.mantisa_a\[8\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
XFILLER_60_266 VPWR VGND sg13g2_decap_8
X_11768_ _05672_ _05669_ _05671_ VPWR VGND sg13g2_nand2_1
X_13507_ VPWR _00058_ net37 VGND sg13g2_inv_1
X_10719_ _04731_ VPWR _04732_ VGND net1821 _04718_ sg13g2_o21ai_1
X_14487_ _00288_ VGND VPWR _01025_ add_result\[12\] clknet_leaf_97_clk sg13g2_dfrbpq_2
X_11699_ _05603_ net1727 _05602_ VPWR VGND sg13g2_nand2_1
XFILLER_127_541 VPWR VGND sg13g2_decap_8
X_13438_ _07098_ net1752 sipo.shift_reg\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_115_725 VPWR VGND sg13g2_decap_8
X_13369_ _07060_ VPWR _00816_ VGND _05357_ net1694 sg13g2_o21ai_1
XFILLER_6_871 VPWR VGND sg13g2_decap_8
XFILLER_114_235 VPWR VGND sg13g2_decap_8
X_07930_ _02205_ fp16_sum_pipe.exp_mant_logic0.b\[10\] VPWR VGND sg13g2_inv_2
XFILLER_87_119 VPWR VGND sg13g2_fill_2
XFILLER_111_964 VPWR VGND sg13g2_decap_8
X_07861_ _02130_ _02048_ _02155_ VPWR VGND sg13g2_nor2_1
XFILLER_96_642 VPWR VGND sg13g2_fill_1
XFILLER_69_878 VPWR VGND sg13g2_decap_8
XFILLER_110_474 VPWR VGND sg13g2_decap_4
X_09600_ VPWR _03717_ _03716_ VGND sg13g2_inv_1
X_07792_ VPWR _02091_ acc_sub.exp_mant_logic0.b\[5\] VGND sg13g2_inv_1
XFILLER_68_388 VPWR VGND sg13g2_fill_1
XFILLER_3_1012 VPWR VGND sg13g2_fill_2
XFILLER_3_1001 VPWR VGND sg13g2_decap_8
XFILLER_110_496 VPWR VGND sg13g2_decap_8
X_09531_ _03648_ _03647_ VPWR VGND sg13g2_inv_2
XFILLER_95_185 VPWR VGND sg13g2_decap_8
XFILLER_52_701 VPWR VGND sg13g2_decap_4
X_09462_ _03592_ VPWR _01254_ VGND net1915 _03591_ sg13g2_o21ai_1
XFILLER_24_425 VPWR VGND sg13g2_fill_1
XFILLER_25_959 VPWR VGND sg13g2_decap_8
X_08413_ _02644_ _02645_ _02647_ _02648_ VPWR VGND sg13g2_nor3_2
X_09393_ _03540_ _03469_ net1738 VPWR VGND sg13g2_nand2_1
X_08344_ _02582_ _02573_ _02587_ _00001_ VPWR VGND sg13g2_nor3_1
XFILLER_33_981 VPWR VGND sg13g2_decap_8
XFILLER_51_299 VPWR VGND sg13g2_decap_8
XFILLER_32_480 VPWR VGND sg13g2_decap_8
X_08275_ _02522_ _02523_ _02524_ VPWR VGND sg13g2_nor2b_1
X_07226_ _01597_ acc_sub.op_sign_logic0.mantisa_a\[0\] acc_sub.op_sign_logic0.mantisa_b\[0\]
+ VPWR VGND sg13g2_nand2_1
X_07157_ _01522_ _01528_ _01529_ VPWR VGND sg13g2_nor2_1
XFILLER_106_758 VPWR VGND sg13g2_decap_8
Xfanout121 net122 net121 VPWR VGND sg13g2_buf_2
Xfanout110 net111 net110 VPWR VGND sg13g2_buf_2
XFILLER_59_300 VPWR VGND sg13g2_decap_8
XFILLER_120_238 VPWR VGND sg13g2_decap_8
Xfanout132 net136 net132 VPWR VGND sg13g2_buf_2
XFILLER_87_653 VPWR VGND sg13g2_fill_2
XFILLER_87_642 VPWR VGND sg13g2_decap_8
XFILLER_47_12 VPWR VGND sg13g2_decap_8
XFILLER_102_986 VPWR VGND sg13g2_decap_8
XFILLER_87_675 VPWR VGND sg13g2_decap_8
XFILLER_86_163 VPWR VGND sg13g2_fill_2
XFILLER_86_152 VPWR VGND sg13g2_decap_8
XFILLER_75_826 VPWR VGND sg13g2_decap_8
XFILLER_59_388 VPWR VGND sg13g2_decap_4
X_09729_ VPWR _03845_ _03844_ VGND sg13g2_inv_1
XFILLER_47_89 VPWR VGND sg13g2_decap_8
XFILLER_90_818 VPWR VGND sg13g2_decap_8
XFILLER_28_786 VPWR VGND sg13g2_fill_2
XFILLER_103_62 VPWR VGND sg13g2_decap_4
X_12740_ _06542_ _06541_ _06513_ VPWR VGND sg13g2_nand2_1
XFILLER_55_594 VPWR VGND sg13g2_decap_4
XFILLER_55_583 VPWR VGND sg13g2_fill_1
XFILLER_15_403 VPWR VGND sg13g2_fill_1
XFILLER_15_414 VPWR VGND sg13g2_fill_2
XFILLER_16_959 VPWR VGND sg13g2_decap_8
X_12671_ VPWR _06485_ div_result\[12\] VGND sg13g2_inv_1
XFILLER_31_907 VPWR VGND sg13g2_decap_8
XFILLER_70_586 VPWR VGND sg13g2_fill_1
XFILLER_63_88 VPWR VGND sg13g2_decap_8
X_14410_ _00211_ VGND VPWR _00949_ fpmul.reg_a_out\[7\] clknet_leaf_127_clk sg13g2_dfrbpq_2
X_11622_ _05527_ _05421_ _05404_ VPWR VGND sg13g2_nand2_1
XFILLER_24_981 VPWR VGND sg13g2_decap_8
X_14341_ _00142_ VGND VPWR _00883_ fpmul.reg_p_out\[5\] clknet_leaf_81_clk sg13g2_dfrbpq_1
XFILLER_8_28 VPWR VGND sg13g2_decap_8
XFILLER_11_653 VPWR VGND sg13g2_decap_4
XFILLER_11_664 VPWR VGND sg13g2_decap_8
XFILLER_11_675 VPWR VGND sg13g2_decap_8
X_11553_ fp16_sum_pipe.add_renorm0.mantisa\[6\] _05427_ fp16_sum_pipe.add_renorm0.mantisa\[7\]
+ _05458_ VPWR VGND sg13g2_a21o_1
X_11484_ _05395_ fp16_res_pipe.x2\[5\] net1945 VPWR VGND sg13g2_nand2_1
X_14272_ _00073_ VGND VPWR _00823_ fp16_res_pipe.x2\[5\] clknet_leaf_18_clk sg13g2_dfrbpq_2
X_10504_ _04548_ _04408_ _04547_ VPWR VGND sg13g2_xnor2_1
XFILLER_6_112 VPWR VGND sg13g2_decap_8
XFILLER_109_552 VPWR VGND sg13g2_fill_2
X_13223_ net3 sipo.bit_counter\[1\] _06949_ _00851_ VPWR VGND sg13g2_a21o_1
X_10435_ _04484_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[4\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[4\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_12_70 VPWR VGND sg13g2_decap_8
X_13154_ _06900_ _06899_ sipo.bit_counter\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_6_189 VPWR VGND sg13g2_fill_2
XFILLER_124_577 VPWR VGND sg13g2_decap_8
XFILLER_112_706 VPWR VGND sg13g2_decap_8
XFILLER_98_918 VPWR VGND sg13g2_decap_8
X_12105_ _05951_ _05949_ _05950_ VPWR VGND sg13g2_nand2_1
X_10366_ _04416_ _04415_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_111_216 VPWR VGND sg13g2_decap_8
X_13085_ _06848_ VPWR _00888_ VGND net1861 _06633_ sg13g2_o21ai_1
XFILLER_3_896 VPWR VGND sg13g2_decap_8
X_10297_ VGND VPWR fp16_res_pipe.exp_mant_logic0.b\[1\] _04177_ _04365_ _04364_ sg13g2_a21oi_1
XFILLER_120_750 VPWR VGND sg13g2_decap_8
XFILLER_78_653 VPWR VGND sg13g2_fill_2
XFILLER_66_804 VPWR VGND sg13g2_decap_8
X_12036_ _05882_ _05880_ _05881_ VPWR VGND sg13g2_nand2_1
XFILLER_2_395 VPWR VGND sg13g2_decap_8
XFILLER_26_7 VPWR VGND sg13g2_decap_8
XFILLER_93_656 VPWR VGND sg13g2_decap_4
XFILLER_81_807 VPWR VGND sg13g2_decap_8
XFILLER_53_509 VPWR VGND sg13g2_decap_8
X_13987_ VPWR _00538_ net9 VGND sg13g2_inv_1
XFILLER_18_252 VPWR VGND sg13g2_decap_8
X_12938_ _06711_ _06710_ net1962 VPWR VGND sg13g2_nand2_1
XFILLER_61_520 VPWR VGND sg13g2_fill_1
X_12869_ _06648_ _06574_ _00014_ VPWR VGND sg13g2_nand2_1
X_14608_ _00409_ VGND VPWR _01140_ fp16_sum_pipe.exp_mant_logic0.a\[3\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_2
XFILLER_21_428 VPWR VGND sg13g2_fill_1
X_14539_ _00340_ VGND VPWR _01075_ acc_sum.op_sign_logic0.mantisa_b\[2\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
XFILLER_30_962 VPWR VGND sg13g2_decap_8
X_08060_ VPWR _02326_ _02314_ VGND sg13g2_inv_1
Xplace1802 acc_sum.seg_reg1.q\[21\] net1802 VPWR VGND sg13g2_buf_2
XFILLER_127_371 VPWR VGND sg13g2_decap_8
Xplace1813 acc_sum.reg1en.q\[0\] net1813 VPWR VGND sg13g2_buf_2
XFILLER_52_0 VPWR VGND sg13g2_decap_8
Xplace1835 fp16_res_pipe.reg3en.q\[0\] net1835 VPWR VGND sg13g2_buf_2
Xplace1824 net1823 net1824 VPWR VGND sg13g2_buf_2
XFILLER_103_717 VPWR VGND sg13g2_decap_8
Xplace1868 fpmul.reg_b_out\[1\] net1868 VPWR VGND sg13g2_buf_2
Xplace1857 fpmul.reg_a_out\[3\] net1857 VPWR VGND sg13g2_buf_2
Xplace1879 net1877 net1879 VPWR VGND sg13g2_buf_2
Xplace1846 net1845 net1846 VPWR VGND sg13g2_buf_2
X_08962_ acc_sub.add_renorm0.exp\[7\] net1699 _03148_ VPWR VGND sg13g2_nor2_1
XFILLER_124_28 VPWR VGND sg13g2_decap_8
X_08893_ VPWR _03080_ _03070_ VGND sg13g2_inv_1
XFILLER_102_249 VPWR VGND sg13g2_fill_1
XFILLER_69_653 VPWR VGND sg13g2_fill_2
XFILLER_69_642 VPWR VGND sg13g2_decap_8
X_07913_ VPWR _02188_ _02187_ VGND sg13g2_inv_1
XFILLER_111_761 VPWR VGND sg13g2_decap_8
X_07844_ _02139_ _01959_ acc_sub.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_97_984 VPWR VGND sg13g2_decap_8
XFILLER_69_675 VPWR VGND sg13g2_fill_1
XFILLER_57_837 VPWR VGND sg13g2_decap_8
XFILLER_56_303 VPWR VGND sg13g2_decap_8
XFILLER_110_282 VPWR VGND sg13g2_fill_1
XFILLER_110_271 VPWR VGND sg13g2_decap_8
XFILLER_84_645 VPWR VGND sg13g2_decap_4
XFILLER_56_336 VPWR VGND sg13g2_decap_8
X_07775_ _02076_ net1649 net1747 VPWR VGND sg13g2_nand2_1
X_09514_ _03631_ acc_sum.add_renorm0.mantisa\[6\] _03623_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_712 VPWR VGND sg13g2_decap_8
XFILLER_24_222 VPWR VGND sg13g2_fill_1
XFILLER_25_767 VPWR VGND sg13g2_decap_8
X_09445_ VPWR _03582_ fp16_res_pipe.add_renorm0.exp\[3\] VGND sg13g2_inv_1
XFILLER_33_14 VPWR VGND sg13g2_decap_8
X_09376_ _03525_ _03382_ _03524_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_288 VPWR VGND sg13g2_decap_8
X_08327_ state\[1\] _02567_ _02572_ VPWR VGND sg13g2_nor2_1
XFILLER_21_973 VPWR VGND sg13g2_decap_8
XFILLER_32_1006 VPWR VGND sg13g2_decap_8
X_08258_ _02459_ _02345_ _02508_ VPWR VGND sg13g2_nor2_1
XFILLER_125_308 VPWR VGND sg13g2_decap_8
X_07209_ _01530_ _01516_ _01581_ VPWR VGND sg13g2_nor2_1
XFILLER_116_5 VPWR VGND sg13g2_decap_8
XFILLER_106_533 VPWR VGND sg13g2_fill_2
XFILLER_4_649 VPWR VGND sg13g2_decap_4
XFILLER_3_126 VPWR VGND sg13g2_decap_8
X_10220_ _04291_ _04292_ _04290_ _04294_ VPWR VGND _04293_ sg13g2_nand4_1
X_08189_ _02262_ _02349_ _02446_ VPWR VGND sg13g2_nor2_1
XFILLER_79_417 VPWR VGND sg13g2_decap_8
XFILLER_0_800 VPWR VGND sg13g2_decap_8
X_10151_ _04138_ _04122_ _04232_ VPWR VGND sg13g2_nor2_1
X_10082_ _04166_ _04167_ _04164_ _04168_ VPWR VGND sg13g2_nand3_1
XFILLER_88_995 VPWR VGND sg13g2_decap_8
XFILLER_87_472 VPWR VGND sg13g2_decap_8
XFILLER_59_152 VPWR VGND sg13g2_fill_2
XFILLER_58_88 VPWR VGND sg13g2_fill_1
X_13910_ VPWR _00461_ net16 VGND sg13g2_inv_1
XFILLER_0_877 VPWR VGND sg13g2_decap_8
X_14890_ _00691_ VGND VPWR _01410_ acc_sub.op_sign_logic0.mantisa_b\[0\] clknet_leaf_61_clk
+ sg13g2_dfrbpq_1
XFILLER_87_483 VPWR VGND sg13g2_decap_4
XFILLER_74_166 VPWR VGND sg13g2_decap_8
X_13841_ VPWR _00392_ net29 VGND sg13g2_inv_1
XFILLER_74_177 VPWR VGND sg13g2_fill_2
XFILLER_62_339 VPWR VGND sg13g2_decap_8
X_13772_ VPWR _00323_ net38 VGND sg13g2_inv_1
XFILLER_56_870 VPWR VGND sg13g2_fill_2
X_10984_ _04978_ fp16_res_pipe.x2\[12\] net1924 VPWR VGND sg13g2_nand2_1
X_12723_ VPWR _06528_ _06428_ VGND sg13g2_inv_1
XFILLER_43_553 VPWR VGND sg13g2_fill_2
X_12654_ _06470_ _05385_ fpdiv.reg_a_out\[13\] VPWR VGND sg13g2_nand2_1
XFILLER_15_288 VPWR VGND sg13g2_decap_8
X_12585_ net1852 _06400_ _06401_ VPWR VGND sg13g2_nor2_2
X_11605_ _05510_ _05465_ _05459_ VPWR VGND sg13g2_nand2_1
XFILLER_30_269 VPWR VGND sg13g2_fill_1
XFILLER_117_809 VPWR VGND sg13g2_decap_8
X_14324_ _00125_ VGND VPWR _00867_ sipo.word\[12\] clknet_leaf_13_clk sg13g2_dfrbpq_2
XFILLER_8_944 VPWR VGND sg13g2_decap_8
XFILLER_12_995 VPWR VGND sg13g2_decap_8
X_11536_ VPWR _05441_ fp16_sum_pipe.add_renorm0.mantisa\[10\] VGND sg13g2_inv_1
XFILLER_23_91 VPWR VGND sg13g2_decap_8
X_14255_ _00056_ VGND VPWR _00806_ acc_sub.x2\[4\] clknet_leaf_20_clk sg13g2_dfrbpq_2
X_13206_ _06938_ VPWR _00857_ VGND _06937_ net1714 sg13g2_o21ai_1
X_11467_ _05386_ fp16_res_pipe.x2\[13\] net1939 VPWR VGND sg13g2_nand2_1
XFILLER_7_498 VPWR VGND sg13g2_decap_8
X_14186_ VPWR _00737_ net116 VGND sg13g2_inv_1
X_11398_ _05343_ VPWR _01069_ VGND _05342_ net1706 sg13g2_o21ai_1
X_10418_ fp16_sum_pipe.reg2en.q\[0\] VPWR _04467_ VGND _04466_ _04384_ sg13g2_o21ai_1
XFILLER_125_886 VPWR VGND sg13g2_decap_8
X_13137_ VPWR _06888_ _06887_ VGND sg13g2_inv_1
XFILLER_3_660 VPWR VGND sg13g2_decap_8
X_10349_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[7\] _04398_ _04399_ VPWR VGND sg13g2_nor2_1
XFILLER_98_759 VPWR VGND sg13g2_decap_4
X_12019_ _05869_ _05845_ _05836_ VPWR VGND sg13g2_nand2_1
XFILLER_39_826 VPWR VGND sg13g2_decap_8
XFILLER_94_954 VPWR VGND sg13g2_decap_8
XFILLER_93_453 VPWR VGND sg13g2_decap_8
XFILLER_93_442 VPWR VGND sg13g2_decap_4
XFILLER_66_656 VPWR VGND sg13g2_decap_8
XFILLER_53_306 VPWR VGND sg13g2_fill_2
XFILLER_38_358 VPWR VGND sg13g2_decap_8
XFILLER_19_550 VPWR VGND sg13g2_fill_1
X_07560_ VPWR _01874_ _01798_ VGND sg13g2_inv_1
XFILLER_0_84 VPWR VGND sg13g2_decap_8
X_07491_ acc_sub.exp_mant_logic0.a\[7\] _01813_ _01814_ VPWR VGND sg13g2_nor2_1
X_09230_ VPWR _03384_ fp16_res_pipe.op_sign_logic0.mantisa_a\[6\] VGND sg13g2_inv_1
XFILLER_61_394 VPWR VGND sg13g2_fill_2
XFILLER_34_597 VPWR VGND sg13g2_decap_8
XFILLER_21_225 VPWR VGND sg13g2_fill_1
X_09161_ _03330_ VPWR _01293_ VGND net1903 _03329_ sg13g2_o21ai_1
X_09092_ _03275_ _03187_ _03194_ VPWR VGND sg13g2_nand2b_1
X_08112_ _02375_ fp16_sum_pipe.exp_mant_logic0.a\[3\] net1684 fp16_sum_pipe.op_sign_logic0.mantisa_a\[6\]
+ net1776 VPWR VGND sg13g2_a22oi_1
XFILLER_30_781 VPWR VGND sg13g2_fill_1
XFILLER_30_792 VPWR VGND sg13g2_decap_4
XFILLER_119_168 VPWR VGND sg13g2_decap_8
XFILLER_119_28 VPWR VGND sg13g2_decap_8
XFILLER_107_308 VPWR VGND sg13g2_fill_1
X_08043_ _02308_ _02245_ _02309_ VPWR VGND sg13g2_nor2_1
XFILLER_116_842 VPWR VGND sg13g2_decap_8
XFILLER_115_341 VPWR VGND sg13g2_decap_8
Xplace1654 _05141_ net1654 VPWR VGND sg13g2_buf_1
Xplace1643 _04158_ net1643 VPWR VGND sg13g2_buf_2
Xplace1665 _01591_ net1665 VPWR VGND sg13g2_buf_2
XFILLER_103_514 VPWR VGND sg13g2_decap_8
Xplace1687 _01840_ net1687 VPWR VGND sg13g2_buf_2
Xplace1676 _06962_ net1676 VPWR VGND sg13g2_buf_2
X_09994_ VPWR _04082_ _04024_ VGND sg13g2_inv_1
XFILLER_103_558 VPWR VGND sg13g2_decap_8
Xplace1698 _05046_ net1698 VPWR VGND sg13g2_buf_2
X_08945_ VGND VPWR _03131_ _03132_ acc_sub.seg_reg1.q\[21\] _03129_ sg13g2_a21oi_2
XFILLER_28_14 VPWR VGND sg13g2_decap_8
X_08876_ VPWR _03063_ _03041_ VGND sg13g2_inv_1
XFILLER_85_943 VPWR VGND sg13g2_decap_8
X_07827_ _01413_ _02122_ _02123_ VPWR VGND sg13g2_nand2_1
XFILLER_84_464 VPWR VGND sg13g2_decap_4
X_07758_ _02061_ net1747 net1651 net1685 net1794 VPWR VGND sg13g2_a22oi_1
XFILLER_84_475 VPWR VGND sg13g2_fill_1
XFILLER_72_615 VPWR VGND sg13g2_decap_8
XFILLER_44_317 VPWR VGND sg13g2_decap_8
XFILLER_44_35 VPWR VGND sg13g2_decap_8
X_07689_ _01998_ acc_sub.exp_mant_logic0.a\[1\] net1672 acc_sub.op_sign_logic0.mantisa_a\[4\]
+ net1780 VPWR VGND sg13g2_a22oi_1
XFILLER_53_884 VPWR VGND sg13g2_fill_1
XFILLER_53_873 VPWR VGND sg13g2_fill_1
XFILLER_13_704 VPWR VGND sg13g2_fill_2
XFILLER_52_394 VPWR VGND sg13g2_decap_8
XFILLER_52_383 VPWR VGND sg13g2_fill_1
X_09428_ _03570_ VPWR _03571_ VGND _03364_ _03566_ sg13g2_o21ai_1
XFILLER_40_556 VPWR VGND sg13g2_decap_8
XFILLER_9_719 VPWR VGND sg13g2_fill_1
X_09359_ _03510_ _03376_ _03509_ VPWR VGND sg13g2_xnor2_1
X_12370_ _06215_ _06214_ _06216_ VPWR VGND sg13g2_xor2_1
Xclkbuf_5_16__f_clk clknet_4_8_0_clk clknet_5_16__leaf_clk VPWR VGND sg13g2_buf_8
X_11321_ _01079_ _05275_ _05276_ VPWR VGND sg13g2_nand2_1
XFILLER_126_639 VPWR VGND sg13g2_decap_8
XFILLER_125_105 VPWR VGND sg13g2_decap_8
XFILLER_4_413 VPWR VGND sg13g2_decap_8
XFILLER_106_330 VPWR VGND sg13g2_fill_2
X_14040_ VPWR _00591_ net74 VGND sg13g2_inv_1
X_11252_ _05209_ _05215_ _05216_ VPWR VGND sg13g2_nor2_1
XFILLER_69_32 VPWR VGND sg13g2_decap_8
XFILLER_5_969 VPWR VGND sg13g2_decap_8
XFILLER_122_812 VPWR VGND sg13g2_decap_8
X_10203_ _04277_ _04278_ _04276_ _04279_ VPWR VGND sg13g2_nand3_1
XFILLER_79_258 VPWR VGND sg13g2_decap_8
XFILLER_69_87 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
X_10134_ net1827 _04128_ _04195_ _04216_ VPWR VGND sg13g2_nand3_1
XFILLER_122_889 VPWR VGND sg13g2_decap_8
XFILLER_121_377 VPWR VGND sg13g2_decap_8
XFILLER_95_718 VPWR VGND sg13g2_decap_8
XFILLER_121_388 VPWR VGND sg13g2_fill_1
X_14942_ _00743_ VGND VPWR _01462_ acc_sub.exp_mant_logic0.a\[10\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_1
XFILLER_94_228 VPWR VGND sg13g2_fill_2
XFILLER_85_31 VPWR VGND sg13g2_decap_8
X_14873_ _00674_ VGND VPWR net1895 acc_sub.reg1en.q\[0\] clknet_leaf_61_clk sg13g2_dfrbpq_2
XFILLER_87_291 VPWR VGND sg13g2_decap_8
XFILLER_85_75 VPWR VGND sg13g2_decap_4
XFILLER_76_976 VPWR VGND sg13g2_fill_1
XFILLER_36_818 VPWR VGND sg13g2_fill_1
XFILLER_76_998 VPWR VGND sg13g2_decap_8
XFILLER_48_689 VPWR VGND sg13g2_fill_2
XFILLER_35_317 VPWR VGND sg13g2_decap_8
X_13824_ VPWR _00375_ net14 VGND sg13g2_inv_1
XFILLER_29_892 VPWR VGND sg13g2_decap_8
XFILLER_91_968 VPWR VGND sg13g2_decap_8
XFILLER_63_659 VPWR VGND sg13g2_fill_1
XFILLER_62_125 VPWR VGND sg13g2_decap_8
X_13755_ VPWR _00306_ net85 VGND sg13g2_inv_1
XFILLER_62_158 VPWR VGND sg13g2_decap_8
X_10967_ fp16_res_pipe.y\[3\] _04686_ net1835 _01124_ VPWR VGND sg13g2_mux2_1
X_13686_ VPWR _00237_ net61 VGND sg13g2_inv_1
X_10898_ _04908_ _04828_ _04791_ VPWR VGND sg13g2_nand2_1
XFILLER_31_523 VPWR VGND sg13g2_decap_8
XFILLER_31_534 VPWR VGND sg13g2_fill_1
XFILLER_31_545 VPWR VGND sg13g2_fill_2
X_12637_ _06435_ _06452_ _06453_ VPWR VGND sg13g2_nor2_1
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
XFILLER_15_1012 VPWR VGND sg13g2_fill_2
XFILLER_31_578 VPWR VGND sg13g2_fill_1
XFILLER_8_730 VPWR VGND sg13g2_fill_1
XFILLER_12_781 VPWR VGND sg13g2_decap_8
XFILLER_31_589 VPWR VGND sg13g2_fill_1
XFILLER_117_617 VPWR VGND sg13g2_fill_2
X_12568_ _06384_ _05387_ fpdiv.reg_a_out\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_7_240 VPWR VGND sg13g2_decap_8
XFILLER_11_280 VPWR VGND sg13g2_decap_4
XFILLER_11_291 VPWR VGND sg13g2_fill_1
X_12499_ VGND VPWR _06332_ net1871 _00958_ _06333_ sg13g2_a21oi_1
X_14307_ _00108_ VGND VPWR _00851_ sipo.bit_counter\[1\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_8_796 VPWR VGND sg13g2_decap_8
X_11519_ _05424_ _05401_ _05423_ VPWR VGND sg13g2_xnor2_1
XFILLER_116_138 VPWR VGND sg13g2_decap_8
X_14238_ _00039_ VGND VPWR _00789_ instr\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_113_823 VPWR VGND sg13g2_decap_8
X_14169_ VPWR _00720_ net101 VGND sg13g2_inv_1
XFILLER_124_182 VPWR VGND sg13g2_decap_8
XFILLER_112_344 VPWR VGND sg13g2_decap_8
XFILLER_112_322 VPWR VGND sg13g2_fill_1
XFILLER_98_556 VPWR VGND sg13g2_decap_8
XFILLER_98_545 VPWR VGND sg13g2_fill_1
XFILLER_3_490 VPWR VGND sg13g2_decap_8
XFILLER_112_399 VPWR VGND sg13g2_decap_8
X_08730_ _02933_ VPWR _01327_ VGND net1815 _02932_ sg13g2_o21ai_1
XFILLER_94_773 VPWR VGND sg13g2_decap_8
X_08661_ _02879_ VPWR _02880_ VGND net1668 _02877_ sg13g2_o21ai_1
XFILLER_66_453 VPWR VGND sg13g2_fill_1
XFILLER_38_133 VPWR VGND sg13g2_decap_8
XFILLER_15_0 VPWR VGND sg13g2_decap_8
XFILLER_27_818 VPWR VGND sg13g2_decap_8
X_07612_ _01926_ _01869_ _01923_ _01871_ net1792 VPWR VGND sg13g2_a22oi_1
XFILLER_93_283 VPWR VGND sg13g2_decap_8
XFILLER_66_486 VPWR VGND sg13g2_fill_1
XFILLER_54_615 VPWR VGND sg13g2_decap_4
XFILLER_93_294 VPWR VGND sg13g2_fill_1
X_08592_ VPWR _02815_ _02814_ VGND sg13g2_inv_1
XFILLER_82_968 VPWR VGND sg13g2_decap_8
X_07543_ _01860_ _01844_ acc_sub.exp_mant_logic0.b\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_81_478 VPWR VGND sg13g2_decap_8
XFILLER_62_670 VPWR VGND sg13g2_fill_1
X_07474_ _01794_ _01796_ _01797_ VPWR VGND sg13g2_nor2_1
XFILLER_62_681 VPWR VGND sg13g2_fill_2
X_09213_ VPWR _03367_ fp16_res_pipe.seg_reg1.q\[20\] VGND sg13g2_inv_1
XFILLER_14_49 VPWR VGND sg13g2_decap_8
X_09144_ acc_sub.reg3en.q\[0\] acc_sub.y\[5\] _03321_ VPWR VGND sg13g2_nor2_1
XFILLER_108_606 VPWR VGND sg13g2_fill_1
X_09075_ VPWR _03259_ acc_sub.y\[12\] VGND sg13g2_inv_1
XFILLER_107_105 VPWR VGND sg13g2_decap_8
X_08026_ _02292_ _02291_ _02223_ VPWR VGND sg13g2_nand2_1
XFILLER_122_119 VPWR VGND sg13g2_decap_8
XFILLER_115_182 VPWR VGND sg13g2_decap_8
XFILLER_104_856 VPWR VGND sg13g2_decap_4
XFILLER_89_589 VPWR VGND sg13g2_fill_1
XFILLER_89_578 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
X_09977_ _04066_ _04067_ _04065_ _01214_ VPWR VGND sg13g2_nand3_1
X_08928_ _03115_ _03004_ _03010_ _02971_ _03009_ VPWR VGND sg13g2_a22oi_1
XFILLER_58_932 VPWR VGND sg13g2_fill_2
XFILLER_85_751 VPWR VGND sg13g2_fill_1
XFILLER_85_740 VPWR VGND sg13g2_decap_8
XFILLER_58_976 VPWR VGND sg13g2_fill_1
X_08859_ VGND VPWR _03045_ _03046_ net1787 _03019_ sg13g2_a21oi_2
XFILLER_84_261 VPWR VGND sg13g2_decap_4
XFILLER_29_155 VPWR VGND sg13g2_decap_8
XFILLER_72_423 VPWR VGND sg13g2_decap_8
XFILLER_55_56 VPWR VGND sg13g2_fill_1
X_11870_ net1850 add_result\[3\] _05763_ VPWR VGND sg13g2_nor2_1
XFILLER_44_147 VPWR VGND sg13g2_decap_8
XFILLER_26_840 VPWR VGND sg13g2_fill_1
XFILLER_72_489 VPWR VGND sg13g2_decap_4
XFILLER_38_1012 VPWR VGND sg13g2_fill_2
XFILLER_38_1001 VPWR VGND sg13g2_decap_8
XFILLER_26_884 VPWR VGND sg13g2_decap_8
X_10821_ VGND VPWR _04831_ _04785_ _04833_ _04832_ sg13g2_a21oi_1
X_13540_ VPWR _00091_ net90 VGND sg13g2_inv_1
XFILLER_71_22 VPWR VGND sg13g2_fill_1
X_10752_ _04765_ _04681_ _04666_ _04670_ _04675_ VPWR VGND sg13g2_a22oi_1
XFILLER_111_84 VPWR VGND sg13g2_decap_8
X_13471_ VPWR _00022_ net82 VGND sg13g2_inv_1
XFILLER_13_545 VPWR VGND sg13g2_fill_2
X_12422_ _06266_ _06267_ _06268_ VPWR VGND sg13g2_nor2_1
XFILLER_40_375 VPWR VGND sg13g2_decap_8
X_10683_ _04696_ _04694_ _04695_ VPWR VGND sg13g2_nand2_1
XFILLER_127_904 VPWR VGND sg13g2_decap_8
XFILLER_126_425 VPWR VGND sg13g2_decap_4
X_12353_ _06199_ _06169_ _06171_ VPWR VGND sg13g2_nand2_1
XFILLER_5_700 VPWR VGND sg13g2_decap_8
XFILLER_114_609 VPWR VGND sg13g2_fill_1
X_12284_ VGND VPWR _06128_ net1869 _06130_ _06129_ sg13g2_a21oi_1
X_11304_ _05262_ net1697 net1812 VPWR VGND sg13g2_nand2_1
XFILLER_5_766 VPWR VGND sg13g2_fill_2
XFILLER_113_119 VPWR VGND sg13g2_decap_8
X_14023_ VPWR _00574_ net100 VGND sg13g2_inv_1
X_11235_ _05198_ _05199_ _05197_ _05200_ VPWR VGND sg13g2_nand3_1
XFILLER_5_799 VPWR VGND sg13g2_decap_4
XFILLER_20_70 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_fill_1
XFILLER_20_92 VPWR VGND sg13g2_decap_8
XFILLER_110_815 VPWR VGND sg13g2_decap_8
X_11166_ _05134_ _05122_ _05135_ VPWR VGND sg13g2_nor2_1
XFILLER_67_206 VPWR VGND sg13g2_decap_4
XFILLER_96_63 VPWR VGND sg13g2_decap_8
X_11097_ _02955_ _02961_ _02953_ _05068_ VPWR VGND sg13g2_nand3_1
XFILLER_1_983 VPWR VGND sg13g2_decap_8
X_10117_ _04197_ _04199_ _04200_ VPWR VGND sg13g2_nor2b_1
XFILLER_121_196 VPWR VGND sg13g2_decap_8
X_14925_ _00726_ VGND VPWR _01445_ fpdiv.divider0.divisor_reg\[5\] clknet_leaf_75_clk
+ sg13g2_dfrbpq_1
XFILLER_76_740 VPWR VGND sg13g2_decap_8
XFILLER_49_965 VPWR VGND sg13g2_fill_2
X_10048_ _04136_ _04124_ _04135_ VPWR VGND sg13g2_nand2_1
XFILLER_75_261 VPWR VGND sg13g2_fill_1
XFILLER_36_626 VPWR VGND sg13g2_decap_8
XFILLER_64_957 VPWR VGND sg13g2_fill_2
X_14856_ _00657_ VGND VPWR _01380_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[7\] clknet_leaf_114_clk
+ sg13g2_dfrbpq_1
XFILLER_90_264 VPWR VGND sg13g2_decap_4
X_13807_ VPWR _00358_ net81 VGND sg13g2_inv_1
X_14787_ _00588_ VGND VPWR _01311_ acc_sum.exp_mant_logic0.a\[0\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
XFILLER_17_884 VPWR VGND sg13g2_decap_8
XFILLER_23_309 VPWR VGND sg13g2_decap_8
XFILLER_91_1003 VPWR VGND sg13g2_decap_8
X_11999_ _05852_ VPWR _05853_ VGND _05827_ _05828_ sg13g2_o21ai_1
XFILLER_44_692 VPWR VGND sg13g2_decap_8
X_13738_ VPWR _00289_ net63 VGND sg13g2_inv_1
XFILLER_31_320 VPWR VGND sg13g2_decap_8
XFILLER_32_865 VPWR VGND sg13g2_fill_1
XFILLER_32_876 VPWR VGND sg13g2_decap_8
X_13669_ VPWR _00220_ net125 VGND sg13g2_inv_1
X_07190_ VPWR _01562_ acc_sub.op_sign_logic0.mantisa_a\[2\] VGND sg13g2_inv_1
XFILLER_118_915 VPWR VGND sg13g2_decap_8
XFILLER_117_414 VPWR VGND sg13g2_fill_2
XFILLER_8_582 VPWR VGND sg13g2_fill_1
XFILLER_126_981 VPWR VGND sg13g2_decap_8
X_09900_ _03994_ _03996_ _03997_ VPWR VGND sg13g2_nor2_1
XFILLER_101_804 VPWR VGND sg13g2_decap_8
X_09831_ net1769 VPWR _03943_ VGND _03942_ _03813_ sg13g2_o21ai_1
XFILLER_98_342 VPWR VGND sg13g2_decap_8
XFILLER_113_686 VPWR VGND sg13g2_decap_8
X_09762_ _03878_ _03851_ _03661_ VPWR VGND sg13g2_xnor2_1
XFILLER_100_314 VPWR VGND sg13g2_decap_8
X_08713_ net1814 acc_sum.add_renorm0.exp\[6\] _02923_ VPWR VGND sg13g2_nor2_1
X_09693_ _03804_ _03808_ _03809_ VPWR VGND sg13g2_nor2_1
XFILLER_27_626 VPWR VGND sg13g2_decap_8
X_08644_ VPWR _02865_ _02800_ VGND sg13g2_inv_1
X_08575_ _02796_ _02798_ _02799_ VPWR VGND sg13g2_nor2_1
XFILLER_82_798 VPWR VGND sg13g2_fill_2
XFILLER_42_629 VPWR VGND sg13g2_fill_1
X_07526_ net1782 _01840_ _01847_ VPWR VGND sg13g2_nor2_2
XFILLER_35_670 VPWR VGND sg13g2_fill_2
XFILLER_23_843 VPWR VGND sg13g2_fill_1
XFILLER_41_14 VPWR VGND sg13g2_decap_8
XFILLER_22_375 VPWR VGND sg13g2_fill_1
XFILLER_23_898 VPWR VGND sg13g2_decap_8
X_07388_ _01734_ net1893 acc\[10\] VPWR VGND sg13g2_nand2_1
X_09127_ _03307_ acc_sub.add_renorm0.exp\[1\] _03306_ VPWR VGND sg13g2_xnor2_1
XFILLER_108_425 VPWR VGND sg13g2_fill_2
XFILLER_124_907 VPWR VGND sg13g2_decap_8
X_09058_ _03243_ VPWR _01309_ VGND net1801 _03138_ sg13g2_o21ai_1
XFILLER_117_970 VPWR VGND sg13g2_decap_8
X_08009_ _02275_ _02223_ VPWR VGND sg13g2_inv_2
XFILLER_116_480 VPWR VGND sg13g2_decap_8
XFILLER_77_504 VPWR VGND sg13g2_decap_8
X_11020_ acc_sum.exp_mant_logic0.b\[12\] _02939_ _04999_ VPWR VGND sg13g2_nor2_1
XFILLER_103_174 VPWR VGND sg13g2_decap_4
XFILLER_89_386 VPWR VGND sg13g2_fill_1
XFILLER_103_196 VPWR VGND sg13g2_decap_8
XFILLER_66_44 VPWR VGND sg13g2_fill_1
XFILLER_85_581 VPWR VGND sg13g2_decap_8
X_12971_ _06740_ _06739_ fp16_sum_pipe.reg1en.d\[0\] _06741_ VPWR VGND sg13g2_a21o_2
XFILLER_66_88 VPWR VGND sg13g2_decap_8
XFILLER_46_924 VPWR VGND sg13g2_fill_1
XFILLER_46_913 VPWR VGND sg13g2_decap_8
X_14710_ _00511_ VGND VPWR _01238_ acc_sum.y\[13\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_73_743 VPWR VGND sg13g2_decap_8
XFILLER_66_99 VPWR VGND sg13g2_fill_2
X_11922_ _05792_ net1882 fpmul.reg_a_out\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_46_957 VPWR VGND sg13g2_fill_2
XFILLER_17_136 VPWR VGND sg13g2_fill_1
XFILLER_18_637 VPWR VGND sg13g2_fill_2
XFILLER_75_1009 VPWR VGND sg13g2_decap_4
XFILLER_60_404 VPWR VGND sg13g2_decap_4
X_14641_ _00442_ VGND VPWR _01173_ fp16_sum_pipe.seg_reg1.q\[20\] clknet_leaf_120_clk
+ sg13g2_dfrbpq_1
XFILLER_17_169 VPWR VGND sg13g2_fill_1
X_11853_ _05750_ VPWR _05751_ VGND _04593_ _05749_ sg13g2_o21ai_1
XFILLER_33_607 VPWR VGND sg13g2_decap_8
XFILLER_73_798 VPWR VGND sg13g2_decap_8
XFILLER_61_949 VPWR VGND sg13g2_fill_1
X_10804_ fp16_res_pipe.add_renorm0.exp\[6\] net1709 _04816_ VPWR VGND sg13g2_nor2_1
XFILLER_14_832 VPWR VGND sg13g2_fill_1
XFILLER_82_87 VPWR VGND sg13g2_fill_2
XFILLER_82_76 VPWR VGND sg13g2_decap_8
X_11784_ _05687_ _05686_ _05627_ VPWR VGND sg13g2_nand2_1
XFILLER_13_320 VPWR VGND sg13g2_decap_8
XFILLER_13_342 VPWR VGND sg13g2_decap_8
XFILLER_25_191 VPWR VGND sg13g2_fill_1
X_14572_ _00373_ VGND VPWR net1933 fp16_sum_pipe.reg1en.q\[0\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_2
X_13523_ VPWR _00074_ net86 VGND sg13g2_inv_1
XFILLER_40_161 VPWR VGND sg13g2_decap_8
X_10735_ _04746_ _04747_ _04748_ VPWR VGND sg13g2_nor2_2
XFILLER_127_701 VPWR VGND sg13g2_decap_8
X_13454_ _07106_ VPWR _00777_ VGND _06927_ net1754 sg13g2_o21ai_1
X_10666_ _04654_ _04678_ _04679_ VPWR VGND sg13g2_nor2_2
X_12405_ _06251_ _06153_ _06250_ VPWR VGND sg13g2_nand2_1
X_13385_ _07069_ net1693 sipo.word\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_115_907 VPWR VGND sg13g2_decap_8
XFILLER_5_541 VPWR VGND sg13g2_decap_8
X_10597_ _04611_ VPWR _01138_ VGND net1934 _02262_ sg13g2_o21ai_1
XFILLER_127_778 VPWR VGND sg13g2_decap_8
XFILLER_126_266 VPWR VGND sg13g2_decap_8
X_12336_ _06182_ _06107_ _06112_ VPWR VGND sg13g2_nand2_1
XFILLER_56_7 VPWR VGND sg13g2_decap_8
XFILLER_99_139 VPWR VGND sg13g2_decap_8
X_12267_ VPWR _06113_ _06112_ VGND sg13g2_inv_1
X_11218_ _05072_ _05183_ _05184_ VPWR VGND sg13g2_nor2_1
X_12198_ VPWR _06044_ _05999_ VGND sg13g2_inv_1
X_14006_ VPWR _00557_ net19 VGND sg13g2_inv_1
XFILLER_123_995 VPWR VGND sg13g2_decap_8
XFILLER_110_601 VPWR VGND sg13g2_decap_4
XFILLER_95_312 VPWR VGND sg13g2_decap_8
X_11149_ _05118_ _05017_ _05119_ VPWR VGND sg13g2_xor2_1
XFILLER_110_656 VPWR VGND sg13g2_decap_8
XFILLER_49_751 VPWR VGND sg13g2_decap_8
XFILLER_76_570 VPWR VGND sg13g2_fill_1
XFILLER_49_773 VPWR VGND sg13g2_decap_8
XFILLER_37_924 VPWR VGND sg13g2_decap_8
XFILLER_36_401 VPWR VGND sg13g2_decap_8
X_14908_ _00709_ VGND VPWR _01428_ acc_sub.op_sign_logic0.mantisa_a\[7\] clknet_leaf_67_clk
+ sg13g2_dfrbpq_1
XFILLER_64_732 VPWR VGND sg13g2_decap_8
XFILLER_48_294 VPWR VGND sg13g2_fill_2
XFILLER_64_787 VPWR VGND sg13g2_fill_2
XFILLER_36_467 VPWR VGND sg13g2_fill_2
X_14839_ _00640_ VGND VPWR _01363_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[1\] clknet_leaf_115_clk
+ sg13g2_dfrbpq_2
X_08360_ _02600_ _02602_ _02599_ _02603_ VPWR VGND sg13g2_nand3_1
XFILLER_51_415 VPWR VGND sg13g2_decap_8
XFILLER_45_990 VPWR VGND sg13g2_decap_8
XFILLER_24_629 VPWR VGND sg13g2_decap_8
X_07311_ _01676_ net1744 _01675_ acc_sub.add_renorm0.mantisa\[5\] net1784 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_60_960 VPWR VGND sg13g2_decap_8
XFILLER_51_459 VPWR VGND sg13g2_decap_8
XFILLER_32_640 VPWR VGND sg13g2_fill_1
X_08291_ _02539_ _02538_ net1638 VPWR VGND sg13g2_nand2_1
X_07242_ _01612_ VPWR _01613_ VGND _01503_ _01505_ sg13g2_o21ai_1
XFILLER_82_0 VPWR VGND sg13g2_decap_4
XFILLER_31_172 VPWR VGND sg13g2_decap_8
XFILLER_118_712 VPWR VGND sg13g2_decap_8
X_07173_ VPWR _01545_ acc_sub.op_sign_logic0.mantisa_b\[0\] VGND sg13g2_inv_1
XFILLER_11_28 VPWR VGND sg13g2_decap_8
XFILLER_127_28 VPWR VGND sg13g2_decap_8
XFILLER_118_789 VPWR VGND sg13g2_decap_8
XFILLER_117_266 VPWR VGND sg13g2_decap_8
XFILLER_106_929 VPWR VGND sg13g2_decap_8
XFILLER_105_406 VPWR VGND sg13g2_decap_8
XFILLER_114_951 VPWR VGND sg13g2_decap_8
X_09814_ net1664 VPWR _03927_ VGND _03916_ _03926_ sg13g2_o21ai_1
XFILLER_100_100 VPWR VGND sg13g2_decap_8
XFILLER_101_667 VPWR VGND sg13g2_decap_4
X_09745_ VPWR _03861_ _03860_ VGND sg13g2_inv_1
XFILLER_101_678 VPWR VGND sg13g2_decap_8
XFILLER_98_1009 VPWR VGND sg13g2_decap_4
XFILLER_28_924 VPWR VGND sg13g2_decap_8
X_09676_ _03792_ _03791_ acc_sum.add_renorm0.exp\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_55_721 VPWR VGND sg13g2_fill_1
XFILLER_36_14 VPWR VGND sg13g2_decap_8
X_08627_ VPWR _02849_ _02848_ VGND sg13g2_inv_1
XFILLER_27_445 VPWR VGND sg13g2_decap_8
XFILLER_54_286 VPWR VGND sg13g2_decap_4
XFILLER_42_437 VPWR VGND sg13g2_decap_8
XFILLER_36_990 VPWR VGND sg13g2_decap_8
XFILLER_27_489 VPWR VGND sg13g2_fill_1
X_08558_ _02775_ _02781_ _02782_ VPWR VGND sg13g2_nor2_1
XFILLER_42_448 VPWR VGND sg13g2_decap_4
X_08489_ _02716_ VPWR _02717_ VGND fpdiv.divider0.remainder_reg\[5\] _02692_ sg13g2_o21ai_1
X_07509_ VGND VPWR _01829_ _01830_ _01831_ _01803_ sg13g2_a21oi_1
XFILLER_52_35 VPWR VGND sg13g2_fill_1
XFILLER_10_301 VPWR VGND sg13g2_decap_8
XFILLER_23_684 VPWR VGND sg13g2_decap_8
X_10520_ VGND VPWR _04560_ net1848 _01165_ _04561_ sg13g2_a21oi_1
XFILLER_23_695 VPWR VGND sg13g2_fill_2
XFILLER_109_723 VPWR VGND sg13g2_fill_1
XFILLER_109_701 VPWR VGND sg13g2_fill_1
XFILLER_108_200 VPWR VGND sg13g2_decap_8
XFILLER_7_839 VPWR VGND sg13g2_decap_8
XFILLER_10_345 VPWR VGND sg13g2_fill_2
XFILLER_11_868 VPWR VGND sg13g2_decap_8
X_10451_ VPWR _04499_ _04468_ VGND sg13g2_inv_1
XFILLER_123_203 VPWR VGND sg13g2_decap_8
X_13170_ VPWR _06914_ sipo.shift_reg\[14\] VGND sg13g2_inv_1
X_10382_ VPWR _04432_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[4\] VGND sg13g2_inv_1
X_12121_ _05967_ net1857 net1866 VPWR VGND sg13g2_nand2_1
XFILLER_2_500 VPWR VGND sg13g2_decap_8
XFILLER_105_951 VPWR VGND sg13g2_decap_8
XFILLER_104_450 VPWR VGND sg13g2_decap_8
XFILLER_81_1013 VPWR VGND sg13g2_fill_1
X_12052_ _05898_ _05889_ _05897_ VPWR VGND sg13g2_nand2_1
XFILLER_120_932 VPWR VGND sg13g2_decap_8
XFILLER_104_461 VPWR VGND sg13g2_fill_1
XFILLER_78_824 VPWR VGND sg13g2_decap_4
X_11003_ _04987_ VPWR _01108_ VGND net1929 _02467_ sg13g2_o21ai_1
XFILLER_93_816 VPWR VGND sg13g2_fill_1
XFILLER_92_315 VPWR VGND sg13g2_decap_8
XFILLER_93_42 VPWR VGND sg13g2_fill_1
X_12954_ _06724_ _06725_ _06715_ _00896_ VPWR VGND sg13g2_nand3_1
XFILLER_58_581 VPWR VGND sg13g2_fill_1
XFILLER_46_743 VPWR VGND sg13g2_fill_2
XFILLER_19_957 VPWR VGND sg13g2_decap_8
XFILLER_73_540 VPWR VGND sg13g2_decap_8
X_11905_ fpmul.seg_reg0.q\[45\] net1854 net1880 _00999_ VPWR VGND sg13g2_mux2_1
XFILLER_46_787 VPWR VGND sg13g2_decap_8
XFILLER_46_754 VPWR VGND sg13g2_fill_2
XFILLER_34_905 VPWR VGND sg13g2_decap_8
X_12885_ acc\[7\] net1907 net1767 _06662_ VPWR VGND sg13g2_nand3_1
XFILLER_45_286 VPWR VGND sg13g2_decap_4
XFILLER_60_245 VPWR VGND sg13g2_decap_8
XFILLER_26_91 VPWR VGND sg13g2_fill_2
X_11836_ _05735_ _05618_ _05617_ VPWR VGND sg13g2_nand2_1
X_14624_ _00425_ VGND VPWR _01156_ fp16_sum_pipe.add_renorm0.exp\[3\] clknet_leaf_120_clk
+ sg13g2_dfrbpq_1
X_14555_ _00356_ VGND VPWR _01091_ acc_sum.op_sign_logic0.mantisa_a\[7\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
XFILLER_42_971 VPWR VGND sg13g2_decap_8
X_11767_ _05670_ VPWR _05671_ VGND net1839 _04585_ sg13g2_o21ai_1
XFILLER_13_150 VPWR VGND sg13g2_fill_2
X_13506_ VPWR _00057_ net37 VGND sg13g2_inv_1
X_10718_ _04731_ _04730_ net1822 VPWR VGND sg13g2_nand2_1
X_14486_ _00287_ VGND VPWR _01024_ add_result\[11\] clknet_leaf_97_clk sg13g2_dfrbpq_2
X_11698_ _05602_ _04587_ _05577_ VPWR VGND sg13g2_xnor2_1
XFILLER_127_520 VPWR VGND sg13g2_decap_8
X_10649_ _04661_ _04650_ _04662_ VPWR VGND sg13g2_and2_1
XFILLER_115_704 VPWR VGND sg13g2_decap_8
X_13368_ _07060_ net1694 sipo.word\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_6_850 VPWR VGND sg13g2_decap_8
XFILLER_127_597 VPWR VGND sg13g2_decap_8
XFILLER_114_214 VPWR VGND sg13g2_decap_8
X_12319_ _06165_ net1860 net1866 VPWR VGND sg13g2_nand2_2
X_13299_ VPWR VGND acc_sub.y\[3\] _07011_ net1711 net1728 _07012_ acc_sum.y\[3\] sg13g2_a221oi_1
XFILLER_5_393 VPWR VGND sg13g2_decap_8
XFILLER_123_792 VPWR VGND sg13g2_decap_8
XFILLER_122_291 VPWR VGND sg13g2_fill_1
XFILLER_122_280 VPWR VGND sg13g2_decap_8
XFILLER_111_943 VPWR VGND sg13g2_decap_8
X_07860_ _02089_ _02015_ _02154_ VPWR VGND sg13g2_nor2_1
X_07791_ _02089_ _01979_ _02090_ VPWR VGND sg13g2_nor2_1
XFILLER_68_367 VPWR VGND sg13g2_decap_8
XFILLER_3_84 VPWR VGND sg13g2_decap_8
X_09530_ _03630_ _03646_ _03647_ VPWR VGND sg13g2_nor2_2
XFILLER_64_551 VPWR VGND sg13g2_decap_4
X_09461_ _03592_ acc_sub.x2\[13\] net1915 VPWR VGND sg13g2_nand2_1
XFILLER_36_242 VPWR VGND sg13g2_fill_2
XFILLER_92_893 VPWR VGND sg13g2_decap_8
XFILLER_92_882 VPWR VGND sg13g2_fill_2
XFILLER_18_990 VPWR VGND sg13g2_decap_8
XFILLER_24_404 VPWR VGND sg13g2_decap_8
XFILLER_25_938 VPWR VGND sg13g2_decap_8
X_08412_ VPWR _02647_ _02646_ VGND sg13g2_inv_1
XFILLER_91_392 VPWR VGND sg13g2_decap_8
X_09392_ VPWR _03539_ _03468_ VGND sg13g2_inv_1
X_08343_ _02582_ _02576_ _02587_ _00000_ VPWR VGND sg13g2_nor3_1
XFILLER_51_278 VPWR VGND sg13g2_decap_8
XFILLER_51_256 VPWR VGND sg13g2_decap_4
XFILLER_33_960 VPWR VGND sg13g2_decap_8
X_08274_ _02523_ _02275_ fp16_sum_pipe.exp_mant_logic0.b\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_20_610 VPWR VGND sg13g2_fill_1
XFILLER_20_632 VPWR VGND sg13g2_fill_1
X_07225_ _01596_ VPWR _01488_ VGND net1798 _01498_ sg13g2_o21ai_1
XFILLER_20_654 VPWR VGND sg13g2_fill_1
XFILLER_22_49 VPWR VGND sg13g2_decap_8
XFILLER_20_687 VPWR VGND sg13g2_fill_2
X_07156_ VPWR _01528_ _01527_ VGND sg13g2_inv_1
XFILLER_121_718 VPWR VGND sg13g2_fill_2
XFILLER_120_217 VPWR VGND sg13g2_decap_8
Xfanout100 net107 net100 VPWR VGND sg13g2_buf_2
XFILLER_87_621 VPWR VGND sg13g2_decap_8
Xfanout122 net128 net122 VPWR VGND sg13g2_buf_2
Xfanout111 net113 net111 VPWR VGND sg13g2_buf_2
Xfanout133 net136 net133 VPWR VGND sg13g2_buf_1
XFILLER_102_965 VPWR VGND sg13g2_decap_8
XFILLER_59_334 VPWR VGND sg13g2_decap_4
XFILLER_74_304 VPWR VGND sg13g2_decap_8
X_09728_ _03844_ _02932_ _03828_ VPWR VGND sg13g2_xnor2_1
XFILLER_86_197 VPWR VGND sg13g2_decap_8
XFILLER_68_890 VPWR VGND sg13g2_decap_8
XFILLER_47_68 VPWR VGND sg13g2_decap_8
X_07989_ _02257_ VPWR _01385_ VGND _02227_ _02248_ sg13g2_o21ai_1
XFILLER_27_231 VPWR VGND sg13g2_fill_2
XFILLER_103_85 VPWR VGND sg13g2_decap_8
X_09659_ _03776_ _03700_ _03711_ VPWR VGND sg13g2_xnor2_1
XFILLER_16_938 VPWR VGND sg13g2_decap_8
XFILLER_103_96 VPWR VGND sg13g2_fill_2
X_12670_ _06484_ VPWR _00939_ VGND _06481_ _06483_ sg13g2_o21ai_1
XFILLER_63_45 VPWR VGND sg13g2_fill_1
XFILLER_43_757 VPWR VGND sg13g2_decap_8
XFILLER_27_297 VPWR VGND sg13g2_decap_8
XFILLER_43_779 VPWR VGND sg13g2_decap_8
X_11621_ VPWR _05526_ _05525_ VGND sg13g2_inv_1
XFILLER_24_960 VPWR VGND sg13g2_decap_8
XFILLER_30_418 VPWR VGND sg13g2_decap_8
X_14340_ _00141_ VGND VPWR _00882_ fpmul.reg_p_out\[4\] clknet_leaf_80_clk sg13g2_dfrbpq_1
XFILLER_23_481 VPWR VGND sg13g2_decap_4
X_11552_ _05450_ _05455_ _05457_ VPWR VGND sg13g2_nor2_2
X_11483_ _05394_ VPWR _01035_ VGND net1948 _05393_ sg13g2_o21ai_1
X_14271_ _00072_ VGND VPWR _00822_ fp16_res_pipe.x2\[4\] clknet_leaf_22_clk sg13g2_dfrbpq_2
X_10503_ _04547_ _04545_ _04546_ _04488_ net1736 VPWR VGND sg13g2_a22oi_1
XFILLER_10_164 VPWR VGND sg13g2_decap_8
X_13222_ _06948_ _06903_ _06945_ _06949_ VPWR VGND sg13g2_nor3_1
XFILLER_6_168 VPWR VGND sg13g2_decap_8
X_10434_ _04482_ VPWR _04483_ VGND _04428_ _04481_ sg13g2_o21ai_1
X_13153_ _06897_ _06898_ _06899_ VPWR VGND sg13g2_nor2_1
X_10365_ VPWR _04415_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[1\] VGND sg13g2_inv_1
X_12104_ _05895_ _05894_ _05892_ _05950_ VPWR VGND sg13g2_nand3_1
XFILLER_97_418 VPWR VGND sg13g2_decap_8
XFILLER_78_610 VPWR VGND sg13g2_fill_2
X_13084_ _06848_ _06847_ _06811_ VPWR VGND sg13g2_nand2_1
XFILLER_3_875 VPWR VGND sg13g2_decap_8
XFILLER_2_374 VPWR VGND sg13g2_decap_8
X_10296_ _04322_ _04233_ _04364_ VPWR VGND sg13g2_nor2_1
XFILLER_78_632 VPWR VGND sg13g2_fill_2
X_12035_ VPWR _05881_ fpmul.reg_a_out\[1\] VGND sg13g2_inv_1
XFILLER_65_304 VPWR VGND sg13g2_fill_2
XFILLER_92_123 VPWR VGND sg13g2_fill_1
XFILLER_19_7 VPWR VGND sg13g2_decap_8
XFILLER_19_721 VPWR VGND sg13g2_fill_1
XFILLER_74_860 VPWR VGND sg13g2_decap_4
X_13986_ VPWR _00537_ net28 VGND sg13g2_inv_1
X_12937_ VPWR _06710_ fpmul.reg_p_out\[3\] VGND sg13g2_inv_1
XFILLER_18_275 VPWR VGND sg13g2_fill_1
XFILLER_19_787 VPWR VGND sg13g2_fill_1
X_12868_ _06647_ _06646_ net1732 VPWR VGND sg13g2_nand2_1
X_11819_ VGND VPWR net1758 _05718_ _05719_ _05572_ sg13g2_a21oi_1
XFILLER_22_919 VPWR VGND sg13g2_decap_8
X_14607_ _00408_ VGND VPWR _01139_ fp16_sum_pipe.exp_mant_logic0.a\[2\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_2
XFILLER_33_267 VPWR VGND sg13g2_decap_4
X_12799_ _06583_ net1910 fp16_res_pipe.y\[14\] VPWR VGND sg13g2_nand2_1
XFILLER_30_941 VPWR VGND sg13g2_decap_8
XFILLER_119_328 VPWR VGND sg13g2_decap_8
X_14538_ _00339_ VGND VPWR _01074_ acc_sum.op_sign_logic0.mantisa_b\[1\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
X_14469_ _00270_ VGND VPWR _01008_ fpmul.result\[15\] clknet_leaf_92_clk sg13g2_dfrbpq_1
XFILLER_127_350 VPWR VGND sg13g2_decap_8
Xplace1803 net1802 net1803 VPWR VGND sg13g2_buf_2
Xplace1814 acc_sum.reg2en.q\[0\] net1814 VPWR VGND sg13g2_buf_1
Xplace1836 fp16_sum_pipe.seg_reg1.q\[21\] net1836 VPWR VGND sg13g2_buf_2
Xplace1825 net1824 net1825 VPWR VGND sg13g2_buf_2
Xplace1869 fpmul.reg_b_out\[0\] net1869 VPWR VGND sg13g2_buf_2
Xplace1858 fpmul.reg_a_out\[2\] net1858 VPWR VGND sg13g2_buf_2
XFILLER_45_0 VPWR VGND sg13g2_decap_8
Xplace1847 fp16_sum_pipe.reg2en.q\[0\] net1847 VPWR VGND sg13g2_buf_2
XFILLER_88_429 VPWR VGND sg13g2_fill_1
XFILLER_88_418 VPWR VGND sg13g2_decap_8
X_08892_ _03075_ _03077_ _03078_ _03079_ VPWR VGND sg13g2_nor3_1
XFILLER_111_740 VPWR VGND sg13g2_decap_8
XFILLER_97_963 VPWR VGND sg13g2_decap_8
X_07912_ fp16_sum_pipe.exp_mant_logic0.b\[13\] _02186_ _02187_ VPWR VGND sg13g2_nor2_1
X_07843_ _01412_ _02137_ _02138_ VPWR VGND sg13g2_nand2_1
XFILLER_112_1006 VPWR VGND sg13g2_decap_8
XFILLER_84_635 VPWR VGND sg13g2_decap_4
XFILLER_68_175 VPWR VGND sg13g2_decap_8
X_07774_ _02075_ net1646 net1794 VPWR VGND sg13g2_nand2_1
XFILLER_84_679 VPWR VGND sg13g2_decap_8
XFILLER_84_668 VPWR VGND sg13g2_fill_1
XFILLER_83_145 VPWR VGND sg13g2_fill_2
X_09513_ _03628_ _03630_ VPWR VGND sg13g2_inv_4
XFILLER_65_882 VPWR VGND sg13g2_decap_8
XFILLER_64_370 VPWR VGND sg13g2_decap_8
XFILLER_17_49 VPWR VGND sg13g2_decap_8
XFILLER_92_690 VPWR VGND sg13g2_decap_4
XFILLER_80_852 VPWR VGND sg13g2_decap_4
XFILLER_80_830 VPWR VGND sg13g2_fill_1
XFILLER_64_392 VPWR VGND sg13g2_fill_1
XFILLER_25_746 VPWR VGND sg13g2_decap_8
X_09444_ _03581_ VPWR _01261_ VGND net1832 _03580_ sg13g2_o21ai_1
XFILLER_52_587 VPWR VGND sg13g2_decap_8
XFILLER_40_727 VPWR VGND sg13g2_fill_2
XFILLER_13_919 VPWR VGND sg13g2_decap_8
XFILLER_40_749 VPWR VGND sg13g2_fill_1
X_09375_ _03523_ VPWR _03524_ VGND net1674 _03521_ sg13g2_o21ai_1
X_08326_ state\[2\] _02559_ _02571_ VPWR VGND sg13g2_nor2_2
XFILLER_20_440 VPWR VGND sg13g2_decap_8
XFILLER_21_952 VPWR VGND sg13g2_decap_8
XFILLER_123_7 VPWR VGND sg13g2_decap_8
X_08257_ _02466_ _02380_ _02507_ VPWR VGND sg13g2_nor2_1
XFILLER_119_884 VPWR VGND sg13g2_decap_8
X_07208_ _01579_ VPWR _01580_ VGND _01516_ _01578_ sg13g2_o21ai_1
X_08188_ _02260_ _02334_ _02445_ VPWR VGND sg13g2_nor2_1
X_07139_ _01511_ _01509_ acc_sub.op_sign_logic0.mantisa_b\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_3_105 VPWR VGND sg13g2_decap_8
X_10150_ _04226_ _04230_ _04231_ VPWR VGND sg13g2_nor2_1
XFILLER_121_537 VPWR VGND sg13g2_fill_2
XFILLER_0_856 VPWR VGND sg13g2_decap_8
X_10081_ _04167_ _04126_ net1828 VPWR VGND sg13g2_nand2_1
XFILLER_88_974 VPWR VGND sg13g2_decap_8
XFILLER_48_849 VPWR VGND sg13g2_decap_8
XFILLER_114_84 VPWR VGND sg13g2_decap_8
XFILLER_101_294 VPWR VGND sg13g2_fill_1
X_13840_ VPWR _00391_ net36 VGND sg13g2_inv_1
XFILLER_74_44 VPWR VGND sg13g2_decap_8
X_13771_ VPWR _00322_ net108 VGND sg13g2_inv_1
XFILLER_16_713 VPWR VGND sg13g2_decap_8
X_10983_ _04977_ VPWR _01118_ VGND net1925 _02464_ sg13g2_o21ai_1
XFILLER_28_584 VPWR VGND sg13g2_fill_1
X_12722_ VPWR _06527_ div_result\[3\] VGND sg13g2_inv_1
XFILLER_43_532 VPWR VGND sg13g2_decap_8
XFILLER_16_735 VPWR VGND sg13g2_decap_8
XFILLER_28_595 VPWR VGND sg13g2_fill_1
XFILLER_90_43 VPWR VGND sg13g2_decap_4
X_12653_ _06408_ _06414_ _06469_ VPWR VGND sg13g2_nor2_1
X_12584_ _06400_ fpdiv.reg_a_out\[7\] fpdiv.reg_b_out\[7\] VPWR VGND sg13g2_xnor2_1
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_11_440 VPWR VGND sg13g2_fill_2
XFILLER_12_974 VPWR VGND sg13g2_decap_8
X_11604_ _05509_ _05483_ _05434_ VPWR VGND sg13g2_nand2_1
X_14323_ _00124_ VGND VPWR _00866_ sipo.word\[11\] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_7_433 VPWR VGND sg13g2_decap_8
X_11535_ fp16_sum_pipe.add_renorm0.mantisa\[9\] _05439_ _05438_ _05440_ VPWR VGND
+ sg13g2_nand3_1
XFILLER_23_70 VPWR VGND sg13g2_decap_8
X_14254_ _00055_ VGND VPWR _00805_ acc_sub.x2\[3\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_11_495 VPWR VGND sg13g2_decap_8
XFILLER_99_52 VPWR VGND sg13g2_fill_2
X_11466_ VPWR _05385_ fpdiv.reg_b_out\[13\] VGND sg13g2_inv_1
X_13205_ _06938_ net1714 sipo.word\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_7_477 VPWR VGND sg13g2_decap_8
XFILLER_125_865 VPWR VGND sg13g2_decap_8
XFILLER_99_85 VPWR VGND sg13g2_fill_2
X_14185_ VPWR _00736_ net116 VGND sg13g2_inv_1
X_11397_ _05343_ net1707 fpdiv.div_out\[8\] VPWR VGND sg13g2_nand2_1
X_10417_ _04466_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[10\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[10\]
+ VPWR VGND sg13g2_nand2_1
X_13136_ _06569_ _06882_ _06887_ VPWR VGND sg13g2_nor2b_1
X_10348_ VPWR _04398_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[7\] VGND sg13g2_inv_1
XFILLER_79_952 VPWR VGND sg13g2_fill_2
X_13067_ fpmul.reg2en.q\[0\] _06834_ _06828_ _06835_ VPWR VGND sg13g2_nand3_1
XFILLER_2_182 VPWR VGND sg13g2_decap_8
X_10279_ _01193_ _04347_ _04348_ VPWR VGND sg13g2_nand2_1
X_12018_ VPWR _05868_ fpmul.seg_reg0.q\[19\] VGND sg13g2_inv_1
XFILLER_39_805 VPWR VGND sg13g2_decap_8
XFILLER_120_570 VPWR VGND sg13g2_fill_1
XFILLER_94_933 VPWR VGND sg13g2_decap_8
XFILLER_93_421 VPWR VGND sg13g2_decap_8
XFILLER_66_635 VPWR VGND sg13g2_decap_8
XFILLER_66_624 VPWR VGND sg13g2_decap_4
XFILLER_65_145 VPWR VGND sg13g2_decap_8
XFILLER_54_819 VPWR VGND sg13g2_decap_8
XFILLER_80_104 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_139_clk clknet_5_2__leaf_clk clknet_leaf_139_clk VPWR VGND sg13g2_buf_8
X_13969_ VPWR _00520_ net18 VGND sg13g2_inv_1
X_07490_ VPWR _01813_ acc_sub.exp_mant_logic0.b\[7\] VGND sg13g2_inv_1
XFILLER_46_381 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_62_885 VPWR VGND sg13g2_decap_8
XFILLER_22_705 VPWR VGND sg13g2_decap_8
X_09160_ _03330_ acc_sub.x2\[14\] net1903 VPWR VGND sg13g2_nand2_1
X_09091_ _03089_ VPWR _03274_ VGND _03262_ _03273_ sg13g2_o21ai_1
X_08111_ _02374_ net1639 _02373_ VPWR VGND sg13g2_nand2_1
XFILLER_119_147 VPWR VGND sg13g2_decap_8
X_08042_ VGND VPWR _02279_ _02230_ _02308_ _02209_ sg13g2_a21oi_1
XFILLER_116_821 VPWR VGND sg13g2_decap_8
XFILLER_115_320 VPWR VGND sg13g2_decap_8
Xplace1644 _04126_ net1644 VPWR VGND sg13g2_buf_1
Xplace1666 net1665 net1666 VPWR VGND sg13g2_buf_1
XFILLER_116_898 VPWR VGND sg13g2_decap_8
XFILLER_115_353 VPWR VGND sg13g2_decap_8
Xplace1677 _06962_ net1677 VPWR VGND sg13g2_buf_1
Xplace1655 _05136_ net1655 VPWR VGND sg13g2_buf_2
X_09993_ VPWR _04081_ _04080_ VGND sg13g2_inv_1
X_08944_ acc_sub.seg_reg1.q\[21\] _03130_ _03036_ _03131_ VPWR VGND sg13g2_nor3_1
Xplace1699 _03146_ net1699 VPWR VGND sg13g2_buf_2
XFILLER_0_119 VPWR VGND sg13g2_decap_8
Xplace1688 _04076_ net1688 VPWR VGND sg13g2_buf_2
XFILLER_88_259 VPWR VGND sg13g2_decap_8
X_08875_ net1790 acc_sub.add_renorm0.mantisa\[10\] _03062_ VPWR VGND sg13g2_nor2_2
XFILLER_85_922 VPWR VGND sg13g2_decap_8
XFILLER_57_646 VPWR VGND sg13g2_fill_1
XFILLER_56_101 VPWR VGND sg13g2_fill_2
XFILLER_29_337 VPWR VGND sg13g2_fill_1
X_07826_ _02123_ acc_sub.exp_mant_logic0.b\[0\] net1669 acc_sub.op_sign_logic0.mantisa_b\[3\]
+ net1781 VPWR VGND sg13g2_a22oi_1
XFILLER_84_443 VPWR VGND sg13g2_decap_8
XFILLER_45_819 VPWR VGND sg13g2_decap_4
X_07757_ _02060_ VPWR _01420_ VGND acc_sub.reg1en.q\[0\] _01501_ sg13g2_o21ai_1
XFILLER_85_999 VPWR VGND sg13g2_decap_8
XFILLER_84_487 VPWR VGND sg13g2_decap_4
XFILLER_56_189 VPWR VGND sg13g2_decap_8
XFILLER_44_307 VPWR VGND sg13g2_fill_2
XFILLER_72_649 VPWR VGND sg13g2_fill_1
XFILLER_44_14 VPWR VGND sg13g2_decap_8
X_07688_ _01997_ _01996_ net1641 VPWR VGND sg13g2_nand2_1
XFILLER_25_565 VPWR VGND sg13g2_decap_8
X_09427_ VGND VPWR _03569_ _03364_ _03570_ net1770 sg13g2_a21oi_1
X_09358_ _03508_ VPWR _03509_ VGND net1674 _03506_ sg13g2_o21ai_1
XFILLER_12_259 VPWR VGND sg13g2_decap_8
XFILLER_100_75 VPWR VGND sg13g2_fill_1
XFILLER_60_35 VPWR VGND sg13g2_decap_8
X_08309_ _02555_ fp16_sum_pipe.exp_mant_logic0.b\[1\] net1658 fp16_sum_pipe.exp_mant_logic0.b\[0\]
+ _02343_ VPWR VGND sg13g2_a22oi_1
XFILLER_126_618 VPWR VGND sg13g2_fill_1
X_11320_ _05276_ acc_sum.exp_mant_logic0.b\[3\] net1681 acc_sum.op_sign_logic0.mantisa_b\[6\]
+ net1762 VPWR VGND sg13g2_a22oi_1
X_09289_ _03443_ _03415_ _03413_ VPWR VGND sg13g2_nand2_2
XFILLER_5_948 VPWR VGND sg13g2_decap_8
XFILLER_107_865 VPWR VGND sg13g2_decap_8
X_11251_ _05215_ _05213_ _05214_ VPWR VGND sg13g2_nand2_1
XFILLER_106_375 VPWR VGND sg13g2_decap_8
X_11182_ _05050_ _05150_ _05151_ VPWR VGND sg13g2_nor2_1
XFILLER_4_469 VPWR VGND sg13g2_decap_8
X_10202_ _04278_ net1688 net1830 VPWR VGND sg13g2_nand2_1
XFILLER_122_868 VPWR VGND sg13g2_decap_8
XFILLER_121_312 VPWR VGND sg13g2_fill_1
XFILLER_79_237 VPWR VGND sg13g2_decap_8
XFILLER_69_99 VPWR VGND sg13g2_decap_4
XFILLER_0_620 VPWR VGND sg13g2_decap_8
X_10133_ _04214_ VPWR _04215_ VGND _03609_ _04175_ sg13g2_o21ai_1
X_14941_ _00742_ VGND VPWR _01461_ acc_sub.exp_mant_logic0.a\[9\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
XFILLER_94_218 VPWR VGND sg13g2_fill_2
XFILLER_88_782 VPWR VGND sg13g2_decap_8
XFILLER_0_675 VPWR VGND sg13g2_fill_1
X_10064_ _04152_ net1637 _04127_ VPWR VGND sg13g2_nand2b_1
X_14872_ _00673_ VGND VPWR net1796 acc_sub.reg2en.q\[0\] clknet_leaf_42_clk sg13g2_dfrbpq_2
XFILLER_63_605 VPWR VGND sg13g2_fill_1
XFILLER_91_947 VPWR VGND sg13g2_decap_8
XFILLER_63_616 VPWR VGND sg13g2_decap_4
X_13823_ VPWR _00374_ net40 VGND sg13g2_inv_1
XFILLER_18_70 VPWR VGND sg13g2_decap_4
XFILLER_44_830 VPWR VGND sg13g2_fill_1
XFILLER_16_510 VPWR VGND sg13g2_fill_1
XFILLER_16_521 VPWR VGND sg13g2_decap_8
X_13754_ VPWR _00305_ net59 VGND sg13g2_inv_1
X_10966_ fp16_res_pipe.y\[4\] _04702_ net1835 _01125_ VPWR VGND sg13g2_mux2_1
XFILLER_16_554 VPWR VGND sg13g2_fill_2
X_12705_ VGND VPWR _06481_ _06513_ _06490_ net1735 sg13g2_a21oi_2
X_13685_ VPWR _00236_ net61 VGND sg13g2_inv_1
X_10897_ VGND VPWR _04906_ _04884_ _04907_ _04774_ sg13g2_a21oi_1
X_12636_ VPWR _06452_ _06451_ VGND sg13g2_inv_1
XFILLER_34_91 VPWR VGND sg13g2_decap_8
XFILLER_86_7 VPWR VGND sg13g2_fill_2
XFILLER_12_760 VPWR VGND sg13g2_decap_8
X_12567_ VGND VPWR _06378_ _06381_ _06383_ _06382_ sg13g2_a21oi_1
X_14306_ _00107_ VGND VPWR _00850_ sipo.bit_counter\[0\] clknet_leaf_9_clk sg13g2_dfrbpq_1
XFILLER_8_753 VPWR VGND sg13g2_decap_4
XFILLER_116_117 VPWR VGND sg13g2_decap_8
X_12498_ net1871 fpmul.seg_reg0.q\[4\] _06333_ VPWR VGND sg13g2_nor2_1
X_11518_ _05423_ _05418_ _05421_ VPWR VGND sg13g2_nand2_1
X_11449_ _05375_ VPWR _01050_ VGND net1947 _05374_ sg13g2_o21ai_1
X_14237_ _00038_ VGND VPWR _00788_ instr\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_124_161 VPWR VGND sg13g2_decap_8
XFILLER_113_802 VPWR VGND sg13g2_decap_8
X_14168_ VPWR _00719_ net103 VGND sg13g2_inv_1
X_13119_ _06874_ VPWR _00880_ VGND net1862 _06721_ sg13g2_o21ai_1
XFILLER_113_879 VPWR VGND sg13g2_decap_8
XFILLER_85_207 VPWR VGND sg13g2_fill_1
XFILLER_39_602 VPWR VGND sg13g2_decap_8
X_14099_ VPWR _00650_ net42 VGND sg13g2_inv_1
XFILLER_85_218 VPWR VGND sg13g2_decap_8
XFILLER_67_933 VPWR VGND sg13g2_decap_8
XFILLER_67_922 VPWR VGND sg13g2_decap_8
XFILLER_39_635 VPWR VGND sg13g2_decap_4
XFILLER_38_112 VPWR VGND sg13g2_decap_8
XFILLER_94_752 VPWR VGND sg13g2_decap_8
X_08660_ _02879_ net1668 _02878_ VPWR VGND sg13g2_nand2_1
XFILLER_94_796 VPWR VGND sg13g2_decap_8
XFILLER_93_262 VPWR VGND sg13g2_decap_8
XFILLER_82_947 VPWR VGND sg13g2_decap_8
XFILLER_81_402 VPWR VGND sg13g2_decap_4
XFILLER_66_465 VPWR VGND sg13g2_decap_8
XFILLER_38_178 VPWR VGND sg13g2_fill_2
X_08591_ _02814_ acc_sum.op_sign_logic0.mantisa_a\[6\] acc_sum.op_sign_logic0.mantisa_b\[6\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_81_446 VPWR VGND sg13g2_decap_8
X_07542_ _01858_ _01859_ _01857_ _01434_ VPWR VGND sg13g2_nand3_1
Xclkbuf_5_22__f_clk clknet_4_11_0_clk clknet_5_22__leaf_clk VPWR VGND sg13g2_buf_8
X_07473_ acc_sub.exp_mant_logic0.a\[12\] _01795_ _01796_ VPWR VGND sg13g2_nor2_1
XFILLER_62_693 VPWR VGND sg13g2_decap_8
XFILLER_61_170 VPWR VGND sg13g2_fill_1
XFILLER_61_192 VPWR VGND sg13g2_fill_1
XFILLER_14_28 VPWR VGND sg13g2_decap_8
X_09212_ VGND VPWR _03359_ _03361_ _01278_ _03365_ sg13g2_a21oi_1
X_09143_ _03320_ VPWR _01301_ VGND net1773 _03113_ sg13g2_o21ai_1
X_09074_ _03258_ VPWR _01308_ VGND net1801 _03244_ sg13g2_o21ai_1
X_08025_ _02291_ _02188_ _02290_ fp16_sum_pipe.exp_mant_logic0.b\[14\] _02238_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_30_49 VPWR VGND sg13g2_decap_8
XFILLER_115_161 VPWR VGND sg13g2_decap_8
XFILLER_103_334 VPWR VGND sg13g2_fill_1
XFILLER_103_312 VPWR VGND sg13g2_decap_8
XFILLER_103_301 VPWR VGND sg13g2_fill_1
XFILLER_39_14 VPWR VGND sg13g2_decap_8
X_09976_ _04067_ net1765 fp16_res_pipe.seg_reg0.q\[23\] VPWR VGND sg13g2_nand2_1
X_08927_ _03114_ _03038_ _03035_ VPWR VGND sg13g2_xnor2_1
X_08858_ net1787 _03044_ _03045_ VPWR VGND sg13g2_nor2_1
XFILLER_84_240 VPWR VGND sg13g2_decap_8
XFILLER_57_454 VPWR VGND sg13g2_decap_8
XFILLER_29_134 VPWR VGND sg13g2_fill_2
X_07809_ _02107_ net1794 _01975_ net1685 acc_sub.exp_mant_logic0.b\[1\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_85_774 VPWR VGND sg13g2_fill_1
XFILLER_73_925 VPWR VGND sg13g2_decap_8
XFILLER_55_35 VPWR VGND sg13g2_decap_8
XFILLER_45_605 VPWR VGND sg13g2_decap_4
X_08789_ _02975_ _02970_ _02976_ VPWR VGND sg13g2_nor2_1
XFILLER_84_295 VPWR VGND sg13g2_fill_2
XFILLER_44_126 VPWR VGND sg13g2_decap_8
XFILLER_38_690 VPWR VGND sg13g2_decap_8
XFILLER_26_863 VPWR VGND sg13g2_decap_8
X_10820_ _04743_ VPWR _04832_ VGND _04785_ _04831_ sg13g2_o21ai_1
XFILLER_125_1005 VPWR VGND sg13g2_decap_8
XFILLER_111_63 VPWR VGND sg13g2_decap_8
X_10751_ _04764_ _04647_ _04679_ _04662_ net1710 VPWR VGND sg13g2_a22oi_1
XFILLER_13_502 VPWR VGND sg13g2_fill_1
X_13470_ VPWR _00021_ net83 VGND sg13g2_inv_1
XFILLER_13_568 VPWR VGND sg13g2_fill_2
X_12421_ VPWR _06267_ _06254_ VGND sg13g2_inv_1
XFILLER_13_579 VPWR VGND sg13g2_fill_1
X_10682_ _04695_ _04642_ VPWR VGND sg13g2_inv_2
X_12352_ _06195_ _06197_ _06198_ VPWR VGND sg13g2_nor2b_1
XFILLER_112_0 VPWR VGND sg13g2_decap_8
XFILLER_107_640 VPWR VGND sg13g2_fill_2
X_12283_ _06089_ _06092_ _06129_ VPWR VGND sg13g2_nor2_1
X_11303_ _05261_ _05124_ net1811 VPWR VGND sg13g2_nand2_1
XFILLER_4_233 VPWR VGND sg13g2_fill_1
X_14022_ VPWR _00573_ net101 VGND sg13g2_inv_1
X_11234_ _05199_ net1810 _05141_ _05075_ acc_sum.exp_mant_logic0.a\[1\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_106_172 VPWR VGND sg13g2_fill_2
XFILLER_96_42 VPWR VGND sg13g2_decap_8
X_11165_ _05134_ _05023_ _05019_ VPWR VGND sg13g2_nand2_1
XFILLER_1_962 VPWR VGND sg13g2_decap_8
XFILLER_122_698 VPWR VGND sg13g2_decap_4
XFILLER_121_175 VPWR VGND sg13g2_decap_8
X_11096_ _05067_ VPWR _01095_ VGND _03343_ _05050_ sg13g2_o21ai_1
X_10116_ VGND VPWR _04177_ net1828 _04199_ _04198_ sg13g2_a21oi_1
X_14924_ _00725_ VGND VPWR _01444_ fpdiv.divider0.divisor_reg\[4\] clknet_leaf_74_clk
+ sg13g2_dfrbpq_1
XFILLER_48_421 VPWR VGND sg13g2_decap_8
X_10047_ _04135_ _04105_ _04134_ VPWR VGND sg13g2_nand2_1
XFILLER_63_402 VPWR VGND sg13g2_decap_8
XFILLER_49_988 VPWR VGND sg13g2_decap_8
XFILLER_90_232 VPWR VGND sg13g2_decap_8
XFILLER_63_424 VPWR VGND sg13g2_fill_1
X_14855_ _00656_ VGND VPWR _01379_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[6\] clknet_leaf_114_clk
+ sg13g2_dfrbpq_1
X_14786_ _00587_ VGND VPWR _01310_ acc_sub.y\[15\] clknet_leaf_39_clk sg13g2_dfrbpq_1
X_13806_ VPWR _00357_ net73 VGND sg13g2_inv_1
X_11998_ _05852_ _05850_ _05851_ VPWR VGND sg13g2_nand2_1
XFILLER_17_863 VPWR VGND sg13g2_decap_8
XFILLER_90_287 VPWR VGND sg13g2_fill_1
XFILLER_72_991 VPWR VGND sg13g2_decap_4
XFILLER_44_682 VPWR VGND sg13g2_decap_8
X_13737_ VPWR _00288_ net55 VGND sg13g2_inv_1
X_10949_ VPWR _04955_ _04748_ VGND sg13g2_inv_1
XFILLER_32_811 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_70_clk clknet_5_30__leaf_clk clknet_leaf_70_clk VPWR VGND sg13g2_buf_8
XFILLER_71_490 VPWR VGND sg13g2_decap_8
X_13668_ VPWR _00219_ net38 VGND sg13g2_inv_1
XFILLER_31_387 VPWR VGND sg13g2_fill_1
X_12619_ _06434_ VPWR _06435_ VGND net1851 fpdiv.div_out\[8\] sg13g2_o21ai_1
X_13599_ VPWR _00150_ net62 VGND sg13g2_inv_1
XFILLER_126_960 VPWR VGND sg13g2_decap_8
XFILLER_6_84 VPWR VGND sg13g2_decap_8
XFILLER_116_19 VPWR VGND sg13g2_decap_8
XFILLER_99_855 VPWR VGND sg13g2_decap_4
X_09830_ _03812_ _03809_ _03942_ VPWR VGND sg13g2_nor2_1
XFILLER_99_866 VPWR VGND sg13g2_decap_8
X_09761_ VPWR _03877_ _03661_ VGND sg13g2_inv_1
XFILLER_101_849 VPWR VGND sg13g2_decap_8
XFILLER_6_1011 VPWR VGND sg13g2_fill_2
X_08712_ VPWR _02922_ acc_sum.seg_reg0.q\[28\] VGND sg13g2_inv_1
XFILLER_79_590 VPWR VGND sg13g2_fill_1
XFILLER_67_741 VPWR VGND sg13g2_fill_2
XFILLER_39_432 VPWR VGND sg13g2_decap_4
XFILLER_39_421 VPWR VGND sg13g2_fill_1
X_09692_ acc_sum.add_renorm0.exp\[1\] _03807_ _03734_ _03808_ VPWR VGND sg13g2_nand3_1
XFILLER_66_251 VPWR VGND sg13g2_decap_8
XFILLER_39_454 VPWR VGND sg13g2_decap_8
X_08643_ VGND VPWR _02854_ _02790_ _02864_ _02789_ sg13g2_a21oi_1
XFILLER_82_733 VPWR VGND sg13g2_decap_8
XFILLER_81_210 VPWR VGND sg13g2_fill_2
XFILLER_26_115 VPWR VGND sg13g2_fill_1
X_08574_ acc_sum.op_sign_logic0.mantisa_a\[10\] _02797_ _02798_ VPWR VGND sg13g2_nor2_2
XFILLER_82_766 VPWR VGND sg13g2_fill_2
XFILLER_81_232 VPWR VGND sg13g2_fill_1
XFILLER_26_159 VPWR VGND sg13g2_fill_2
X_07525_ _01846_ _01844_ acc_sub.exp_mant_logic0.b\[12\] VPWR VGND sg13g2_nand2_1
XFILLER_34_170 VPWR VGND sg13g2_decap_8
XFILLER_22_310 VPWR VGND sg13g2_decap_8
XFILLER_25_49 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_61_clk clknet_5_28__leaf_clk clknet_leaf_61_clk VPWR VGND sg13g2_buf_8
X_07456_ acc_sub.reg1en.q\[0\] _01779_ VPWR VGND sg13g2_inv_4
XFILLER_50_674 VPWR VGND sg13g2_fill_2
XFILLER_50_663 VPWR VGND sg13g2_decap_8
XFILLER_23_877 VPWR VGND sg13g2_decap_8
X_07387_ VPWR _01733_ acc_sub.exp_mant_logic0.a\[10\] VGND sg13g2_inv_1
XFILLER_6_509 VPWR VGND sg13g2_decap_8
XFILLER_10_538 VPWR VGND sg13g2_decap_4
X_09126_ VGND VPWR _03080_ _03225_ _03306_ _03224_ sg13g2_a21oi_1
XFILLER_109_949 VPWR VGND sg13g2_decap_8
XFILLER_108_404 VPWR VGND sg13g2_decap_8
X_09057_ _03243_ _03215_ _03242_ VPWR VGND sg13g2_nand2_1
XFILLER_108_448 VPWR VGND sg13g2_decap_4
XFILLER_123_407 VPWR VGND sg13g2_decap_4
X_08008_ _02274_ VPWR _01383_ VGND fp16_sum_pipe.reg1en.q\[0\] _02259_ sg13g2_o21ai_1
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_89_365 VPWR VGND sg13g2_fill_1
XFILLER_89_354 VPWR VGND sg13g2_decap_8
XFILLER_1_258 VPWR VGND sg13g2_fill_1
XFILLER_104_687 VPWR VGND sg13g2_decap_4
X_09959_ _04052_ _04054_ VPWR VGND sg13g2_inv_4
XFILLER_92_508 VPWR VGND sg13g2_fill_1
XFILLER_73_700 VPWR VGND sg13g2_decap_8
XFILLER_66_67 VPWR VGND sg13g2_decap_8
XFILLER_66_56 VPWR VGND sg13g2_fill_2
XFILLER_58_763 VPWR VGND sg13g2_fill_2
XFILLER_57_240 VPWR VGND sg13g2_decap_8
X_12970_ _06740_ net1910 fp16_res_pipe.y\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_18_627 VPWR VGND sg13g2_fill_1
XFILLER_58_796 VPWR VGND sg13g2_fill_1
XFILLER_45_446 VPWR VGND sg13g2_decap_8
X_11921_ VPWR _05791_ fpmul.seg_reg0.q\[39\] VGND sg13g2_inv_1
XFILLER_61_917 VPWR VGND sg13g2_decap_4
XFILLER_17_159 VPWR VGND sg13g2_fill_2
X_14640_ _00441_ VGND VPWR _01172_ fp16_sum_pipe.add_renorm0.mantisa\[11\] clknet_leaf_110_clk
+ sg13g2_dfrbpq_2
X_11852_ VGND VPWR _05749_ _04593_ _05750_ fp16_sum_pipe.seg_reg1.q\[21\] sg13g2_a21oi_1
XFILLER_122_84 VPWR VGND sg13g2_decap_8
XFILLER_61_939 VPWR VGND sg13g2_fill_1
X_14571_ _00372_ VGND VPWR net1843 fp16_sum_pipe.reg2en.q\[0\] clknet_leaf_120_clk
+ sg13g2_dfrbpq_2
X_10803_ VPWR _04815_ _04814_ VGND sg13g2_inv_1
Xclkbuf_leaf_52_clk clknet_5_19__leaf_clk clknet_leaf_52_clk VPWR VGND sg13g2_buf_8
X_13522_ VPWR _00073_ net84 VGND sg13g2_inv_1
X_11783_ VPWR _05686_ _05624_ VGND sg13g2_inv_1
XFILLER_41_674 VPWR VGND sg13g2_decap_8
XFILLER_40_140 VPWR VGND sg13g2_decap_8
XFILLER_14_888 VPWR VGND sg13g2_decap_8
X_10734_ VPWR _04747_ _04717_ VGND sg13g2_inv_1
X_13453_ _07106_ net1754 sipo.shift_reg\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_9_336 VPWR VGND sg13g2_decap_8
XFILLER_9_358 VPWR VGND sg13g2_decap_8
X_10665_ VPWR _04678_ _04658_ VGND sg13g2_inv_1
XFILLER_13_387 VPWR VGND sg13g2_decap_8
X_12404_ _06247_ _06249_ _06250_ VPWR VGND sg13g2_nor2b_2
X_13384_ _07068_ VPWR _00809_ VGND _03603_ net1695 sg13g2_o21ai_1
XFILLER_9_369 VPWR VGND sg13g2_fill_1
XFILLER_127_757 VPWR VGND sg13g2_decap_8
X_12335_ VGND VPWR _06174_ _06177_ _06181_ _06180_ sg13g2_a21oi_1
XFILLER_5_520 VPWR VGND sg13g2_decap_8
XFILLER_31_70 VPWR VGND sg13g2_decap_8
X_10596_ _04611_ acc_sub.x2\[1\] net1933 VPWR VGND sg13g2_nand2_1
XFILLER_126_245 VPWR VGND sg13g2_decap_8
XFILLER_31_81 VPWR VGND sg13g2_fill_2
XFILLER_108_993 VPWR VGND sg13g2_decap_8
X_12266_ _06104_ _06105_ _06088_ _06112_ VPWR VGND sg13g2_nand3_1
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_5_575 VPWR VGND sg13g2_fill_2
XFILLER_123_974 VPWR VGND sg13g2_decap_8
X_11217_ VPWR _05183_ _05181_ VGND sg13g2_inv_1
X_12197_ _06043_ _06041_ _06042_ VPWR VGND sg13g2_nand2_1
X_14005_ VPWR _00556_ net19 VGND sg13g2_inv_1
XFILLER_122_484 VPWR VGND sg13g2_decap_8
XFILLER_110_624 VPWR VGND sg13g2_fill_1
X_11148_ _05117_ VPWR _05118_ VGND _05030_ net1698 sg13g2_o21ai_1
X_11079_ _05055_ VPWR _01100_ VGND _03333_ _05050_ sg13g2_o21ai_1
XFILLER_48_251 VPWR VGND sg13g2_decap_8
XFILLER_37_903 VPWR VGND sg13g2_decap_8
X_14907_ _00708_ VGND VPWR _01427_ acc_sub.op_sign_logic0.mantisa_a\[6\] clknet_leaf_68_clk
+ sg13g2_dfrbpq_2
XFILLER_36_446 VPWR VGND sg13g2_decap_8
X_14838_ _00639_ VGND VPWR _01362_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[0\] clknet_leaf_116_clk
+ sg13g2_dfrbpq_1
XFILLER_63_265 VPWR VGND sg13g2_fill_2
X_07310_ _01675_ _01535_ _01605_ VPWR VGND sg13g2_xnor2_1
XFILLER_108_1000 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_43_clk clknet_5_23__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
X_14769_ _00570_ VGND VPWR _01293_ acc_sum.exp_mant_logic0.b\[14\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_2
X_08290_ _02534_ _02537_ _02533_ _02538_ VPWR VGND sg13g2_nand3_1
X_07241_ _01612_ _01611_ _01508_ VPWR VGND sg13g2_nand2_1
XFILLER_20_847 VPWR VGND sg13g2_fill_2
X_07172_ VPWR _01544_ _01543_ VGND sg13g2_inv_1
XFILLER_75_0 VPWR VGND sg13g2_decap_4
XFILLER_118_768 VPWR VGND sg13g2_decap_8
XFILLER_106_908 VPWR VGND sg13g2_decap_8
XFILLER_9_892 VPWR VGND sg13g2_decap_8
XFILLER_117_245 VPWR VGND sg13g2_decap_8
XFILLER_114_930 VPWR VGND sg13g2_decap_8
XFILLER_28_1001 VPWR VGND sg13g2_decap_8
XFILLER_28_1012 VPWR VGND sg13g2_fill_2
XFILLER_113_473 VPWR VGND sg13g2_decap_8
X_09813_ _03908_ _03925_ _03926_ VPWR VGND sg13g2_nor2_1
XFILLER_101_602 VPWR VGND sg13g2_decap_8
XFILLER_99_696 VPWR VGND sg13g2_fill_2
XFILLER_98_162 VPWR VGND sg13g2_decap_8
XFILLER_59_516 VPWR VGND sg13g2_fill_2
XFILLER_101_646 VPWR VGND sg13g2_fill_2
XFILLER_101_635 VPWR VGND sg13g2_decap_8
XFILLER_87_858 VPWR VGND sg13g2_decap_4
XFILLER_86_357 VPWR VGND sg13g2_fill_2
XFILLER_59_549 VPWR VGND sg13g2_decap_4
X_09744_ _03838_ _03859_ _03860_ VPWR VGND sg13g2_nor2_2
XFILLER_100_156 VPWR VGND sg13g2_fill_2
XFILLER_100_145 VPWR VGND sg13g2_decap_8
XFILLER_95_880 VPWR VGND sg13g2_fill_1
XFILLER_86_368 VPWR VGND sg13g2_fill_2
XFILLER_74_519 VPWR VGND sg13g2_decap_8
XFILLER_67_560 VPWR VGND sg13g2_fill_2
XFILLER_55_711 VPWR VGND sg13g2_fill_2
XFILLER_28_903 VPWR VGND sg13g2_decap_8
X_09675_ _02924_ _03790_ _03791_ VPWR VGND sg13g2_nor2_1
XFILLER_54_210 VPWR VGND sg13g2_decap_8
XFILLER_39_284 VPWR VGND sg13g2_decap_8
XFILLER_82_563 VPWR VGND sg13g2_fill_2
X_08626_ VGND VPWR _02847_ _02751_ _02848_ _02750_ sg13g2_a21oi_1
XFILLER_54_243 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_34_clk clknet_5_20__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
X_08557_ VPWR _02781_ _02780_ VGND sg13g2_inv_1
XFILLER_52_14 VPWR VGND sg13g2_decap_8
X_08488_ _02692_ VPWR _02716_ VGND _02665_ _02715_ sg13g2_o21ai_1
X_07508_ VPWR _01830_ _01805_ VGND sg13g2_inv_1
XFILLER_122_1008 VPWR VGND sg13g2_decap_4
X_07439_ VGND VPWR _01768_ net1749 _01447_ _01769_ sg13g2_a21oi_1
XFILLER_10_324 VPWR VGND sg13g2_decap_4
XFILLER_11_847 VPWR VGND sg13g2_decap_8
XFILLER_22_184 VPWR VGND sg13g2_fill_2
XFILLER_7_818 VPWR VGND sg13g2_decap_8
XFILLER_22_195 VPWR VGND sg13g2_fill_2
X_10450_ VGND VPWR _04462_ _04465_ _01172_ _04498_ sg13g2_a21oi_1
X_09109_ _03219_ _03229_ _03291_ VPWR VGND sg13g2_nor2_1
X_10381_ _04430_ VPWR _04431_ VGND _04418_ _04429_ sg13g2_o21ai_1
XFILLER_105_930 VPWR VGND sg13g2_decap_8
X_12120_ _05966_ fpmul.reg_a_out\[6\] net1867 VPWR VGND sg13g2_nand2_1
XFILLER_123_259 VPWR VGND sg13g2_decap_8
X_12051_ VGND VPWR _05892_ _05894_ _05897_ _05896_ sg13g2_a21oi_1
XFILLER_2_556 VPWR VGND sg13g2_decap_8
XFILLER_120_911 VPWR VGND sg13g2_decap_8
XFILLER_117_84 VPWR VGND sg13g2_decap_8
XFILLER_78_847 VPWR VGND sg13g2_decap_8
XFILLER_78_814 VPWR VGND sg13g2_fill_1
XFILLER_77_33 VPWR VGND sg13g2_decap_8
X_11002_ _04987_ fp16_res_pipe.x2\[3\] net1928 VPWR VGND sg13g2_nand2_1
XFILLER_77_324 VPWR VGND sg13g2_fill_2
XFILLER_120_988 VPWR VGND sg13g2_decap_8
X_12953_ _06725_ net1717 _00007_ VPWR VGND sg13g2_nand2_1
XFILLER_18_413 VPWR VGND sg13g2_decap_4
XFILLER_19_936 VPWR VGND sg13g2_decap_8
X_11904_ fpmul.seg_reg0.q\[46\] fpmul.reg_a_out\[7\] net1876 _01000_ VPWR VGND sg13g2_mux2_1
XFILLER_45_232 VPWR VGND sg13g2_decap_4
XFILLER_61_725 VPWR VGND sg13g2_decap_8
X_12884_ VGND VPWR net1936 add_result\[7\] _06661_ net1950 sg13g2_a21oi_1
XFILLER_45_265 VPWR VGND sg13g2_decap_8
X_14623_ _00424_ VGND VPWR _01155_ fp16_sum_pipe.add_renorm0.exp\[2\] clknet_leaf_111_clk
+ sg13g2_dfrbpq_1
XFILLER_33_416 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_5_17__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_26_70 VPWR VGND sg13g2_decap_8
X_11835_ VGND VPWR _05506_ _05598_ _05734_ _05733_ sg13g2_a21oi_1
X_14554_ _00355_ VGND VPWR _01090_ acc_sum.op_sign_logic0.mantisa_a\[6\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_11766_ _05670_ _05606_ net1839 VPWR VGND sg13g2_nand2_1
X_13505_ VPWR _00056_ net82 VGND sg13g2_inv_1
X_14485_ _00286_ VGND VPWR _01023_ add_result\[10\] clknet_leaf_100_clk sg13g2_dfrbpq_2
XFILLER_9_133 VPWR VGND sg13g2_decap_8
X_10717_ _04727_ _04728_ _04721_ _04730_ VPWR VGND _04729_ sg13g2_nand4_1
XFILLER_13_162 VPWR VGND sg13g2_decap_8
X_13436_ _06906_ VPWR _00785_ VGND _06911_ _06905_ sg13g2_o21ai_1
X_11697_ VPWR _05601_ _05599_ VGND sg13g2_inv_1
XFILLER_42_91 VPWR VGND sg13g2_decap_8
X_10648_ fp16_res_pipe.add_renorm0.mantisa\[7\] _04646_ fp16_res_pipe.add_renorm0.mantisa\[8\]
+ _04661_ VPWR VGND sg13g2_a21o_1
XFILLER_9_199 VPWR VGND sg13g2_decap_8
XFILLER_127_576 VPWR VGND sg13g2_decap_8
X_13367_ _07059_ VPWR _00817_ VGND _03327_ net1696 sg13g2_o21ai_1
X_10579_ _04602_ VPWR _01147_ VGND net1930 _02203_ sg13g2_o21ai_1
XFILLER_10_891 VPWR VGND sg13g2_decap_8
X_13298_ _07010_ _06952_ _07011_ VPWR VGND sg13g2_nor2_1
X_12318_ VPWR _06164_ _06163_ VGND sg13g2_inv_1
XFILLER_69_803 VPWR VGND sg13g2_fill_2
X_12249_ _06095_ _05956_ _05962_ VPWR VGND sg13g2_nand2_1
XFILLER_123_771 VPWR VGND sg13g2_decap_8
XFILLER_111_922 VPWR VGND sg13g2_decap_8
XFILLER_69_836 VPWR VGND sg13g2_decap_8
XFILLER_110_421 VPWR VGND sg13g2_fill_1
XFILLER_110_410 VPWR VGND sg13g2_decap_8
XFILLER_3_63 VPWR VGND sg13g2_decap_8
XFILLER_111_999 VPWR VGND sg13g2_decap_8
X_07790_ _02089_ acc_sub.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_inv_2
XFILLER_95_154 VPWR VGND sg13g2_decap_8
XFILLER_84_817 VPWR VGND sg13g2_decap_8
XFILLER_77_891 VPWR VGND sg13g2_fill_2
XFILLER_49_593 VPWR VGND sg13g2_decap_8
XFILLER_64_541 VPWR VGND sg13g2_decap_8
X_09460_ VPWR _03591_ fp16_res_pipe.exp_mant_logic0.a\[13\] VGND sg13g2_inv_1
XFILLER_25_917 VPWR VGND sg13g2_decap_8
X_08411_ fpdiv.divider0.counter\[1\] fpdiv.divider0.counter\[0\] _02646_ VPWR VGND
+ sg13g2_nor2_1
XFILLER_36_254 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_16_clk clknet_5_6__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
XFILLER_51_246 VPWR VGND sg13g2_decap_4
X_09391_ _03537_ VPWR _03538_ VGND _03397_ _03536_ sg13g2_o21ai_1
X_08342_ _02583_ _02584_ _02585_ _02586_ _02587_ VPWR VGND sg13g2_nor4_1
X_08273_ _02466_ _02396_ _02522_ VPWR VGND sg13g2_nor2_1
X_07224_ _01595_ VPWR _01596_ VGND acc_sub.op_sign_logic0.s_a _01591_ sg13g2_o21ai_1
XFILLER_22_28 VPWR VGND sg13g2_decap_8
XFILLER_118_521 VPWR VGND sg13g2_fill_2
X_07155_ _01524_ _01526_ _01527_ VPWR VGND sg13g2_nor2_2
XFILLER_118_576 VPWR VGND sg13g2_decap_8
Xfanout101 net102 net101 VPWR VGND sg13g2_buf_2
Xfanout112 net113 net112 VPWR VGND sg13g2_buf_1
XFILLER_113_281 VPWR VGND sg13g2_fill_2
Xfanout134 net136 net134 VPWR VGND sg13g2_buf_2
XFILLER_102_944 VPWR VGND sg13g2_decap_8
XFILLER_87_655 VPWR VGND sg13g2_fill_1
Xfanout123 net124 net123 VPWR VGND sg13g2_buf_2
XFILLER_101_454 VPWR VGND sg13g2_decap_4
XFILLER_87_666 VPWR VGND sg13g2_decap_4
X_07988_ _02257_ fp16_sum_pipe.exp_mant_logic0.a\[8\] _02250_ fp16_sum_pipe.seg_reg0.q\[23\]
+ net1775 VPWR VGND sg13g2_a22oi_1
X_09727_ _03840_ _03842_ _03843_ VPWR VGND sg13g2_nor2_1
XFILLER_101_498 VPWR VGND sg13g2_decap_8
XFILLER_47_47 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_decap_8
XFILLER_16_917 VPWR VGND sg13g2_decap_8
XFILLER_27_221 VPWR VGND sg13g2_fill_1
X_09658_ VGND VPWR _03774_ _03775_ net1802 _03770_ sg13g2_a21oi_2
XFILLER_103_53 VPWR VGND sg13g2_decap_4
XFILLER_82_371 VPWR VGND sg13g2_fill_2
XFILLER_82_360 VPWR VGND sg13g2_decap_8
XFILLER_43_736 VPWR VGND sg13g2_decap_8
XFILLER_43_725 VPWR VGND sg13g2_decap_8
XFILLER_27_276 VPWR VGND sg13g2_decap_8
XFILLER_28_799 VPWR VGND sg13g2_decap_4
X_09589_ _03705_ VPWR _03706_ VGND net1805 _03650_ sg13g2_o21ai_1
X_08609_ _02832_ _02744_ _02831_ _02815_ _02726_ VPWR VGND sg13g2_a22oi_1
XFILLER_70_555 VPWR VGND sg13g2_fill_2
X_11620_ net1838 fp16_sum_pipe.add_renorm0.mantisa\[10\] _05525_ VPWR VGND sg13g2_nor2_1
XFILLER_51_791 VPWR VGND sg13g2_fill_2
X_10502_ VGND VPWR net1673 _04447_ _04546_ net1736 sg13g2_a21oi_1
X_11482_ _05394_ fp16_res_pipe.x2\[6\] net1948 VPWR VGND sg13g2_nand2_1
X_14270_ _00071_ VGND VPWR _00821_ fp16_res_pipe.x2\[3\] clknet_leaf_20_clk sg13g2_dfrbpq_2
XFILLER_7_626 VPWR VGND sg13g2_fill_2
XFILLER_109_565 VPWR VGND sg13g2_decap_8
X_13221_ sipo.bit_counter\[1\] sipo.bit_counter\[0\] _06948_ VPWR VGND sg13g2_nor2_1
XFILLER_6_147 VPWR VGND sg13g2_decap_8
X_10433_ _04482_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[3\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[3\]
+ VPWR VGND sg13g2_nand2_1
X_13152_ _06898_ sipo.bit_counter\[1\] sipo.bit_counter\[0\] VPWR VGND sg13g2_nand2_1
X_10364_ _04414_ _04413_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_124_557 VPWR VGND sg13g2_decap_4
XFILLER_88_43 VPWR VGND sg13g2_decap_8
X_12103_ _05949_ _05948_ _05893_ VPWR VGND sg13g2_nand2_1
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_3_854 VPWR VGND sg13g2_decap_8
XFILLER_88_98 VPWR VGND sg13g2_decap_8
X_13083_ VGND VPWR _06809_ _06761_ _06847_ _06835_ sg13g2_a21oi_1
XFILLER_2_353 VPWR VGND sg13g2_decap_8
X_10295_ _04361_ _04362_ _04363_ VPWR VGND sg13g2_nor2_1
XFILLER_104_270 VPWR VGND sg13g2_decap_4
XFILLER_78_644 VPWR VGND sg13g2_fill_1
X_12034_ _05880_ fpmul.reg_a_out\[2\] net1863 VPWR VGND sg13g2_nand2_1
XFILLER_93_614 VPWR VGND sg13g2_fill_2
XFILLER_120_785 VPWR VGND sg13g2_decap_8
XFILLER_77_198 VPWR VGND sg13g2_fill_1
XFILLER_77_176 VPWR VGND sg13g2_decap_8
XFILLER_59_891 VPWR VGND sg13g2_decap_8
XFILLER_18_210 VPWR VGND sg13g2_decap_4
XFILLER_58_390 VPWR VGND sg13g2_fill_2
XFILLER_19_744 VPWR VGND sg13g2_decap_8
Xclkbuf_5_3__f_clk clknet_4_1_0_clk clknet_5_3__leaf_clk VPWR VGND sg13g2_buf_8
X_13985_ VPWR _00536_ net28 VGND sg13g2_inv_1
XFILLER_92_179 VPWR VGND sg13g2_fill_1
XFILLER_92_168 VPWR VGND sg13g2_decap_8
XFILLER_80_308 VPWR VGND sg13g2_decap_8
X_12936_ _06709_ _06705_ _06708_ _06527_ net1948 VPWR VGND sg13g2_a22oi_1
XFILLER_74_894 VPWR VGND sg13g2_decap_4
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_19_799 VPWR VGND sg13g2_decap_8
X_12867_ _06645_ VPWR _06646_ VGND net1960 _06643_ sg13g2_o21ai_1
XFILLER_61_533 VPWR VGND sg13g2_decap_8
XFILLER_61_588 VPWR VGND sg13g2_decap_8
X_11818_ _05718_ _05658_ _05667_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_1011 VPWR VGND sg13g2_fill_2
X_14606_ _00407_ VGND VPWR _01138_ fp16_sum_pipe.exp_mant_logic0.a\[1\] clknet_leaf_119_clk
+ sg13g2_dfrbpq_2
XFILLER_33_257 VPWR VGND sg13g2_fill_1
X_14537_ _00338_ VGND VPWR _01073_ acc_sum.op_sign_logic0.mantisa_b\[0\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_2
X_12798_ acc\[14\] net1908 net1767 _06582_ VPWR VGND sg13g2_nand3_1
XFILLER_15_994 VPWR VGND sg13g2_decap_8
XFILLER_30_920 VPWR VGND sg13g2_decap_8
X_11749_ _05653_ _05625_ net1839 VPWR VGND sg13g2_nand2_1
XFILLER_88_1009 VPWR VGND sg13g2_decap_4
X_14468_ _00269_ VGND VPWR _01007_ fpmul.seg_reg0.q\[53\] clknet_leaf_125_clk sg13g2_dfrbpq_1
XFILLER_30_997 VPWR VGND sg13g2_decap_8
X_14399_ _00200_ VGND VPWR _00938_ div_result\[12\] clknet_leaf_89_clk sg13g2_dfrbpq_1
X_13419_ _07088_ VPWR _00794_ VGND _07044_ net1722 sg13g2_o21ai_1
Xplace1804 net1802 net1804 VPWR VGND sg13g2_buf_1
Xplace1815 net1814 net1815 VPWR VGND sg13g2_buf_1
Xplace1826 fp16_res_pipe.add_renorm0.mantisa\[11\] net1826 VPWR VGND sg13g2_buf_2
XFILLER_115_568 VPWR VGND sg13g2_fill_2
XFILLER_89_909 VPWR VGND sg13g2_decap_8
Xplace1859 fpmul.reg_a_out\[1\] net1859 VPWR VGND sg13g2_buf_2
Xplace1848 net1847 net1848 VPWR VGND sg13g2_buf_2
Xplace1837 net1836 net1837 VPWR VGND sg13g2_buf_2
X_08960_ _03146_ _03145_ VPWR VGND sg13g2_inv_2
Xclkbuf_leaf_5_clk clknet_5_5__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_08891_ _03059_ _03076_ _03078_ VPWR VGND sg13g2_nor2_1
XFILLER_97_942 VPWR VGND sg13g2_decap_8
X_07911_ _02186_ fp16_sum_pipe.exp_mant_logic0.a\[13\] VPWR VGND sg13g2_inv_2
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_07842_ _02138_ net1779 acc_sub.op_sign_logic0.mantisa_b\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_110_251 VPWR VGND sg13g2_fill_1
XFILLER_68_154 VPWR VGND sg13g2_decap_8
XFILLER_57_828 VPWR VGND sg13g2_decap_4
XFILLER_111_796 VPWR VGND sg13g2_decap_8
XFILLER_83_124 VPWR VGND sg13g2_decap_8
XFILLER_110_295 VPWR VGND sg13g2_decap_8
X_07773_ _02073_ _01821_ _02074_ VPWR VGND sg13g2_nor2_1
XFILLER_17_28 VPWR VGND sg13g2_decap_8
XFILLER_92_680 VPWR VGND sg13g2_decap_8
X_09443_ _03581_ net1833 fp16_res_pipe.seg_reg0.q\[26\] VPWR VGND sg13g2_nand2_1
XFILLER_80_875 VPWR VGND sg13g2_decap_8
XFILLER_40_706 VPWR VGND sg13g2_decap_8
X_09374_ net1674 VPWR _03523_ VGND _03387_ _03522_ sg13g2_o21ai_1
XFILLER_24_268 VPWR VGND sg13g2_decap_4
XFILLER_71_1013 VPWR VGND sg13g2_fill_1
XFILLER_33_791 VPWR VGND sg13g2_fill_1
XFILLER_21_931 VPWR VGND sg13g2_decap_8
XFILLER_33_49 VPWR VGND sg13g2_decap_8
XFILLER_32_290 VPWR VGND sg13g2_fill_1
X_08256_ _02468_ _02322_ _02506_ VPWR VGND sg13g2_nor2_1
XFILLER_119_863 VPWR VGND sg13g2_decap_8
X_07207_ _01511_ VPWR _01579_ VGND _01510_ _01504_ sg13g2_o21ai_1
X_08187_ _01374_ _02443_ _02444_ VPWR VGND sg13g2_nand2_1
XFILLER_118_373 VPWR VGND sg13g2_decap_8
X_07138_ acc_sub.op_sign_logic0.mantisa_b\[9\] _01509_ _01510_ VPWR VGND sg13g2_nor2_1
XFILLER_106_579 VPWR VGND sg13g2_decap_8
XFILLER_88_953 VPWR VGND sg13g2_decap_8
XFILLER_87_430 VPWR VGND sg13g2_decap_8
XFILLER_59_121 VPWR VGND sg13g2_fill_1
XFILLER_0_835 VPWR VGND sg13g2_decap_8
X_10080_ _04166_ _04165_ net1746 VPWR VGND sg13g2_nand2_1
XFILLER_102_763 VPWR VGND sg13g2_decap_8
XFILLER_59_154 VPWR VGND sg13g2_fill_1
XFILLER_58_57 VPWR VGND sg13g2_fill_2
XFILLER_75_647 VPWR VGND sg13g2_fill_1
XFILLER_114_63 VPWR VGND sg13g2_decap_8
XFILLER_74_23 VPWR VGND sg13g2_decap_8
XFILLER_63_809 VPWR VGND sg13g2_fill_2
XFILLER_74_67 VPWR VGND sg13g2_decap_8
X_13770_ VPWR _00321_ net109 VGND sg13g2_inv_1
XFILLER_62_308 VPWR VGND sg13g2_decap_8
XFILLER_56_894 VPWR VGND sg13g2_fill_1
XFILLER_56_883 VPWR VGND sg13g2_decap_8
X_10982_ _04977_ fp16_res_pipe.x2\[13\] net1925 VPWR VGND sg13g2_nand2_1
X_12721_ _06526_ VPWR _00930_ VGND _06520_ net1741 sg13g2_o21ai_1
X_12652_ _06468_ _06467_ _06415_ VPWR VGND sg13g2_nand2b_1
XFILLER_90_22 VPWR VGND sg13g2_fill_1
XFILLER_43_588 VPWR VGND sg13g2_fill_2
X_11603_ VGND VPWR _05506_ _05470_ _05508_ _05507_ sg13g2_a21oi_1
XFILLER_24_780 VPWR VGND sg13g2_decap_8
XFILLER_24_791 VPWR VGND sg13g2_fill_2
XFILLER_30_205 VPWR VGND sg13g2_decap_8
XFILLER_31_739 VPWR VGND sg13g2_decap_8
X_12583_ _06399_ _06398_ _06378_ VPWR VGND sg13g2_nand2b_1
XFILLER_8_902 VPWR VGND sg13g2_decap_8
XFILLER_12_953 VPWR VGND sg13g2_decap_8
X_14322_ _00123_ VGND VPWR _00865_ sipo.word\[10\] clknet_leaf_13_clk sg13g2_dfrbpq_2
X_11534_ _05439_ _05431_ _05426_ VPWR VGND sg13g2_nand2_1
X_14253_ _00054_ VGND VPWR _00804_ acc_sub.x2\[2\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_11465_ fpdiv.reg_b_out\[14\] fp16_res_pipe.x2\[14\] net1942 _01043_ VPWR VGND sg13g2_mux2_1
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_7_456 VPWR VGND sg13g2_decap_8
XFILLER_99_42 VPWR VGND sg13g2_fill_1
X_13204_ VPWR _06937_ sipo.shift_reg\[3\] VGND sg13g2_inv_1
X_10416_ net1838 _04465_ VPWR VGND sg13g2_inv_4
XFILLER_125_844 VPWR VGND sg13g2_decap_8
XFILLER_124_343 VPWR VGND sg13g2_fill_1
XFILLER_99_97 VPWR VGND sg13g2_decap_4
X_14184_ VPWR _00735_ net116 VGND sg13g2_inv_1
X_11396_ _05342_ fpdiv.div_out\[7\] VPWR VGND sg13g2_inv_2
X_13135_ _06884_ _06886_ _00876_ VPWR VGND sg13g2_nor2_1
X_10347_ _04394_ _04396_ _04397_ VPWR VGND sg13g2_nor2_2
XFILLER_78_430 VPWR VGND sg13g2_decap_8
X_13066_ VPWR _06834_ _06833_ VGND sg13g2_inv_1
XFILLER_2_161 VPWR VGND sg13g2_decap_8
X_10278_ _04348_ net1763 fp16_res_pipe.op_sign_logic0.mantisa_b\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_31_7 VPWR VGND sg13g2_decap_8
XFILLER_94_912 VPWR VGND sg13g2_decap_8
XFILLER_78_452 VPWR VGND sg13g2_fill_1
XFILLER_78_441 VPWR VGND sg13g2_fill_1
XFILLER_66_603 VPWR VGND sg13g2_decap_8
X_12017_ VGND VPWR _05866_ net1877 _00974_ _05867_ sg13g2_a21oi_1
XFILLER_94_989 VPWR VGND sg13g2_decap_8
XFILLER_65_124 VPWR VGND sg13g2_decap_8
XFILLER_65_179 VPWR VGND sg13g2_fill_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_19_563 VPWR VGND sg13g2_decap_8
XFILLER_19_574 VPWR VGND sg13g2_fill_2
X_13968_ VPWR _00519_ net7 VGND sg13g2_inv_1
X_12919_ _00010_ net1731 net1702 _06693_ VPWR VGND sg13g2_nand3_1
XFILLER_62_820 VPWR VGND sg13g2_decap_8
XFILLER_19_596 VPWR VGND sg13g2_fill_2
XFILLER_62_875 VPWR VGND sg13g2_fill_2
XFILLER_61_363 VPWR VGND sg13g2_fill_2
XFILLER_61_341 VPWR VGND sg13g2_decap_8
XFILLER_55_1008 VPWR VGND sg13g2_decap_4
X_13899_ VPWR _00450_ net12 VGND sg13g2_inv_1
XFILLER_15_780 VPWR VGND sg13g2_decap_8
XFILLER_15_791 VPWR VGND sg13g2_fill_1
XFILLER_14_290 VPWR VGND sg13g2_fill_2
X_09090_ _03195_ _03180_ _03273_ VPWR VGND sg13g2_nor2_1
XFILLER_119_126 VPWR VGND sg13g2_decap_8
XFILLER_9_84 VPWR VGND sg13g2_decap_8
X_08110_ _02371_ _02372_ _02370_ _02373_ VPWR VGND sg13g2_nand3_1
X_08041_ _02307_ _02305_ VPWR VGND sg13g2_inv_2
XFILLER_116_800 VPWR VGND sg13g2_decap_8
Xplace1634 _05256_ net1634 VPWR VGND sg13g2_buf_2
Xplace1645 _02324_ net1645 VPWR VGND sg13g2_buf_2
Xplace1667 net1666 net1667 VPWR VGND sg13g2_buf_2
XFILLER_116_877 VPWR VGND sg13g2_decap_8
Xplace1678 net1677 net1678 VPWR VGND sg13g2_buf_2
XFILLER_89_739 VPWR VGND sg13g2_decap_4
Xplace1656 net1655 net1656 VPWR VGND sg13g2_buf_1
X_09992_ _04079_ VPWR _04080_ VGND fp16_res_pipe.exp_mant_logic0.a\[8\] _04034_ sg13g2_o21ai_1
X_08943_ _03034_ _03032_ _03130_ VPWR VGND sg13g2_nor2_1
XFILLER_103_549 VPWR VGND sg13g2_decap_4
Xplace1689 _04050_ net1689 VPWR VGND sg13g2_buf_2
Xclkbuf_4_15_0_clk clknet_0_clk clknet_4_15_0_clk VPWR VGND sg13g2_buf_8
XFILLER_97_772 VPWR VGND sg13g2_decap_8
XFILLER_97_750 VPWR VGND sg13g2_decap_4
X_08874_ _03060_ _03058_ _03061_ VPWR VGND sg13g2_nor2_1
XFILLER_84_422 VPWR VGND sg13g2_decap_8
XFILLER_57_625 VPWR VGND sg13g2_decap_8
XFILLER_57_614 VPWR VGND sg13g2_decap_4
X_07825_ _02122_ _02121_ net1640 VPWR VGND sg13g2_nand2_1
XFILLER_85_978 VPWR VGND sg13g2_decap_8
XFILLER_28_49 VPWR VGND sg13g2_decap_8
X_07756_ net1796 _02058_ net1686 _02060_ VPWR VGND sg13g2_nand3_1
XFILLER_38_883 VPWR VGND sg13g2_decap_8
XFILLER_53_842 VPWR VGND sg13g2_fill_2
XFILLER_25_511 VPWR VGND sg13g2_decap_8
X_07687_ _01994_ _01995_ _01993_ _01996_ VPWR VGND sg13g2_nand3_1
XFILLER_64_190 VPWR VGND sg13g2_decap_8
XFILLER_52_341 VPWR VGND sg13g2_fill_2
X_09426_ _03568_ _03443_ _03569_ VPWR VGND sg13g2_xor2_1
XFILLER_13_706 VPWR VGND sg13g2_fill_1
XFILLER_80_672 VPWR VGND sg13g2_decap_8
XFILLER_40_514 VPWR VGND sg13g2_decap_4
XFILLER_12_216 VPWR VGND sg13g2_decap_4
X_09357_ _03508_ net1674 _03507_ VPWR VGND sg13g2_nand2b_1
X_09288_ _03397_ _03441_ _03408_ _03442_ VPWR VGND sg13g2_nor3_1
X_08308_ _02554_ fp16_sum_pipe.exp_mant_logic0.b\[4\] _02408_ net1842 _02332_ VPWR
+ VGND sg13g2_a22oi_1
XFILLER_20_260 VPWR VGND sg13g2_decap_4
XFILLER_60_69 VPWR VGND sg13g2_decap_8
XFILLER_60_58 VPWR VGND sg13g2_decap_4
X_08239_ _02491_ fp16_sum_pipe.exp_mant_logic0.b\[4\] net1645 _02343_ fp16_sum_pipe.exp_mant_logic0.b\[6\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_119_682 VPWR VGND sg13g2_decap_8
XFILLER_5_927 VPWR VGND sg13g2_decap_8
XFILLER_109_63 VPWR VGND sg13g2_decap_8
XFILLER_107_844 VPWR VGND sg13g2_decap_8
X_11250_ _05214_ net1653 net1809 VPWR VGND sg13g2_nand2_1
XFILLER_4_448 VPWR VGND sg13g2_decap_8
XFILLER_106_354 VPWR VGND sg13g2_decap_8
X_11181_ _05133_ _05149_ _05150_ VPWR VGND sg13g2_nor2_1
X_10201_ _04277_ net1643 net1745 VPWR VGND sg13g2_nand2_1
XFILLER_122_847 VPWR VGND sg13g2_decap_8
XFILLER_79_216 VPWR VGND sg13g2_decap_8
X_10132_ _04214_ net1643 fp16_res_pipe.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_0_665 VPWR VGND sg13g2_decap_4
XFILLER_125_84 VPWR VGND sg13g2_decap_8
X_14940_ _00741_ VGND VPWR _01460_ acc_sub.exp_mant_logic0.a\[8\] clknet_leaf_45_clk
+ sg13g2_dfrbpq_2
XFILLER_85_11 VPWR VGND sg13g2_fill_2
XFILLER_75_422 VPWR VGND sg13g2_decap_8
XFILLER_0_698 VPWR VGND sg13g2_decap_8
X_14871_ _00672_ VGND VPWR net1797 acc_sub.reg3en.q\[0\] clknet_leaf_46_clk sg13g2_dfrbpq_2
XFILLER_75_444 VPWR VGND sg13g2_fill_2
XFILLER_48_647 VPWR VGND sg13g2_decap_4
XFILLER_47_124 VPWR VGND sg13g2_decap_8
XFILLER_36_809 VPWR VGND sg13g2_decap_8
XFILLER_16_500 VPWR VGND sg13g2_decap_4
XFILLER_29_883 VPWR VGND sg13g2_fill_1
X_13822_ VPWR _00373_ net44 VGND sg13g2_inv_1
X_13753_ VPWR _00304_ net59 VGND sg13g2_inv_1
XFILLER_28_382 VPWR VGND sg13g2_decap_8
X_12704_ _06512_ _06456_ _06511_ VPWR VGND sg13g2_xnor2_1
XFILLER_44_875 VPWR VGND sg13g2_decap_8
XFILLER_43_341 VPWR VGND sg13g2_decap_8
X_10965_ fp16_res_pipe.y\[5\] _04768_ fp16_res_pipe.reg3en.q\[0\] _01126_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_16_544 VPWR VGND sg13g2_fill_1
XFILLER_71_694 VPWR VGND sg13g2_decap_8
XFILLER_71_672 VPWR VGND sg13g2_decap_8
X_13684_ VPWR _00235_ net61 VGND sg13g2_inv_1
XFILLER_44_886 VPWR VGND sg13g2_fill_2
XFILLER_43_374 VPWR VGND sg13g2_decap_8
X_10896_ _04791_ VPWR _04906_ VGND _04796_ _04812_ sg13g2_o21ai_1
X_12635_ _06437_ _06450_ _06451_ VPWR VGND sg13g2_nor2_1
XFILLER_70_182 VPWR VGND sg13g2_fill_1
XFILLER_34_70 VPWR VGND sg13g2_decap_8
XFILLER_31_569 VPWR VGND sg13g2_decap_8
X_12566_ _06379_ _06380_ _06382_ VPWR VGND sg13g2_nor2b_1
X_14305_ _00106_ VGND VPWR _00849_ acc\[15\] clknet_leaf_50_clk sg13g2_dfrbpq_2
XFILLER_8_765 VPWR VGND sg13g2_decap_4
XFILLER_117_619 VPWR VGND sg13g2_fill_1
X_12497_ _06332_ _06330_ _06331_ VPWR VGND sg13g2_xnor2_1
X_11448_ _05375_ acc_sub.x2\[5\] net1946 VPWR VGND sg13g2_nand2_1
X_14236_ _00037_ VGND VPWR _00787_ instr\[1\] clknet_leaf_19_clk sg13g2_dfrbpq_2
XFILLER_50_91 VPWR VGND sg13g2_decap_8
XFILLER_125_674 VPWR VGND sg13g2_decap_8
XFILLER_124_140 VPWR VGND sg13g2_decap_8
X_14167_ VPWR _00718_ net90 VGND sg13g2_inv_1
X_11379_ _05330_ net1762 acc_sum.op_sign_logic0.mantisa_b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_113_858 VPWR VGND sg13g2_decap_8
X_13118_ net1700 _06870_ _06802_ _06874_ VPWR VGND _06873_ sg13g2_nand4_1
XFILLER_4_993 VPWR VGND sg13g2_decap_8
XFILLER_79_761 VPWR VGND sg13g2_decap_8
XFILLER_61_1012 VPWR VGND sg13g2_fill_2
X_14098_ VPWR _00649_ net43 VGND sg13g2_inv_1
XFILLER_100_519 VPWR VGND sg13g2_decap_8
XFILLER_79_794 VPWR VGND sg13g2_decap_8
XFILLER_79_772 VPWR VGND sg13g2_fill_2
X_13049_ VPWR _06817_ _06816_ VGND sg13g2_inv_1
XFILLER_93_230 VPWR VGND sg13g2_fill_2
XFILLER_66_444 VPWR VGND sg13g2_decap_8
XFILLER_39_669 VPWR VGND sg13g2_fill_1
XFILLER_39_658 VPWR VGND sg13g2_decap_8
X_08590_ acc_sum.op_sign_logic0.mantisa_a\[7\] acc_sum.op_sign_logic0.mantisa_b\[7\]
+ _02813_ VPWR VGND sg13g2_nor2_1
XFILLER_82_926 VPWR VGND sg13g2_decap_8
X_07541_ _01859_ _01779_ acc_sub.seg_reg0.q\[24\] VPWR VGND sg13g2_nand2_1
XFILLER_66_499 VPWR VGND sg13g2_decap_8
XFILLER_35_831 VPWR VGND sg13g2_fill_1
XFILLER_19_382 VPWR VGND sg13g2_decap_8
XFILLER_53_149 VPWR VGND sg13g2_decap_8
XFILLER_35_875 VPWR VGND sg13g2_decap_4
XFILLER_90_981 VPWR VGND sg13g2_decap_8
X_07472_ VPWR _01795_ acc_sub.exp_mant_logic0.b\[12\] VGND sg13g2_inv_1
XFILLER_35_897 VPWR VGND sg13g2_decap_8
XFILLER_34_385 VPWR VGND sg13g2_fill_2
XFILLER_22_514 VPWR VGND sg13g2_fill_2
X_09142_ _03320_ net1773 acc_sub.y\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_30_580 VPWR VGND sg13g2_decap_8
X_09073_ _03258_ _03255_ _03257_ VPWR VGND sg13g2_nand2_1
XFILLER_30_28 VPWR VGND sg13g2_decap_8
X_08024_ _02290_ _02289_ _02189_ VPWR VGND sg13g2_nand2_1
XFILLER_116_663 VPWR VGND sg13g2_decap_4
XFILLER_115_140 VPWR VGND sg13g2_decap_8
XFILLER_2_919 VPWR VGND sg13g2_decap_8
XFILLER_118_1013 VPWR VGND sg13g2_fill_1
XFILLER_104_847 VPWR VGND sg13g2_decap_4
XFILLER_89_547 VPWR VGND sg13g2_fill_2
XFILLER_1_429 VPWR VGND sg13g2_decap_8
X_09975_ _04066_ _04056_ fp16_res_pipe.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
X_08926_ VGND VPWR _03109_ net1787 _03113_ _03112_ sg13g2_a21oi_1
XFILLER_112_880 VPWR VGND sg13g2_decap_8
XFILLER_58_934 VPWR VGND sg13g2_fill_1
X_08857_ _03044_ _03021_ _03042_ VPWR VGND sg13g2_xnor2_1
XFILLER_111_390 VPWR VGND sg13g2_fill_1
X_07808_ _02106_ acc_sub.exp_mant_logic0.b\[4\] net1649 acc_sub.exp_mant_logic0.b\[2\]
+ net1651 VPWR VGND sg13g2_a22oi_1
XFILLER_85_786 VPWR VGND sg13g2_decap_4
XFILLER_58_989 VPWR VGND sg13g2_fill_2
XFILLER_57_466 VPWR VGND sg13g2_decap_8
XFILLER_55_14 VPWR VGND sg13g2_decap_8
XFILLER_29_168 VPWR VGND sg13g2_decap_4
X_08788_ VPWR _02975_ acc_sub.add_renorm0.mantisa\[6\] VGND sg13g2_inv_1
XFILLER_84_274 VPWR VGND sg13g2_decap_4
XFILLER_73_959 VPWR VGND sg13g2_decap_8
XFILLER_44_105 VPWR VGND sg13g2_decap_8
X_07739_ _02044_ _02018_ net1793 VPWR VGND sg13g2_nand2_1
XFILLER_72_469 VPWR VGND sg13g2_fill_2
XFILLER_72_458 VPWR VGND sg13g2_decap_8
XFILLER_37_190 VPWR VGND sg13g2_fill_1
XFILLER_111_42 VPWR VGND sg13g2_decap_8
XFILLER_81_992 VPWR VGND sg13g2_decap_8
XFILLER_41_834 VPWR VGND sg13g2_fill_2
XFILLER_40_311 VPWR VGND sg13g2_fill_2
X_10750_ _04763_ _04695_ _04720_ _04672_ _04694_ VPWR VGND sg13g2_a22oi_1
XFILLER_25_385 VPWR VGND sg13g2_fill_2
XFILLER_40_344 VPWR VGND sg13g2_fill_1
XFILLER_40_333 VPWR VGND sg13g2_decap_8
XFILLER_40_322 VPWR VGND sg13g2_fill_1
X_09409_ _03553_ VPWR _03554_ VGND _03464_ _03552_ sg13g2_o21ai_1
XFILLER_13_547 VPWR VGND sg13g2_fill_1
X_10681_ net1710 _04693_ _04694_ VPWR VGND sg13g2_nor2_2
XFILLER_71_68 VPWR VGND sg13g2_fill_2
X_12420_ net1854 fpmul.reg_b_out\[6\] _06266_ VPWR VGND sg13g2_nor2_1
XFILLER_127_939 VPWR VGND sg13g2_decap_8
X_12351_ _06197_ _06164_ _06196_ VPWR VGND sg13g2_xnor2_1
X_12282_ _06128_ _06092_ _06089_ VPWR VGND sg13g2_nand2_1
X_11302_ _05260_ net1656 _05253_ VPWR VGND sg13g2_nand2_1
XFILLER_122_600 VPWR VGND sg13g2_decap_4
XFILLER_105_0 VPWR VGND sg13g2_decap_8
X_14021_ VPWR _00572_ net101 VGND sg13g2_inv_1
XFILLER_84_1012 VPWR VGND sg13g2_fill_2
XFILLER_84_1001 VPWR VGND sg13g2_decap_8
X_11233_ _05198_ acc_sum.exp_mant_logic0.a\[2\] _05161_ net1653 net1808 VPWR VGND
+ sg13g2_a22oi_1
XFILLER_122_644 VPWR VGND sg13g2_decap_4
X_11164_ _05133_ _05132_ _05129_ VPWR VGND sg13g2_nand2b_1
XFILLER_68_709 VPWR VGND sg13g2_decap_8
XFILLER_1_941 VPWR VGND sg13g2_decap_8
XFILLER_121_154 VPWR VGND sg13g2_decap_8
X_11095_ _05067_ acc_sum.exp_mant_logic0.a\[7\] _05052_ net1760 acc_sum.seg_reg0.q\[22\]
+ VPWR VGND sg13g2_a22oi_1
X_10115_ _03615_ net1703 _04198_ VPWR VGND sg13g2_nor2_1
X_14923_ _00724_ VGND VPWR _01443_ acc_sub.reg_add_sub.q\[0\] clknet_leaf_61_clk sg13g2_dfrbpq_1
XFILLER_102_390 VPWR VGND sg13g2_decap_4
XFILLER_49_967 VPWR VGND sg13g2_fill_1
XFILLER_49_945 VPWR VGND sg13g2_decap_8
XFILLER_0_484 VPWR VGND sg13g2_decap_8
XFILLER_29_70 VPWR VGND sg13g2_fill_2
X_10046_ _04017_ _04115_ _04119_ _04134_ VPWR VGND sg13g2_nor3_1
XFILLER_91_712 VPWR VGND sg13g2_decap_4
XFILLER_75_252 VPWR VGND sg13g2_decap_8
XFILLER_48_466 VPWR VGND sg13g2_decap_8
XFILLER_36_617 VPWR VGND sg13g2_decap_4
XFILLER_36_606 VPWR VGND sg13g2_decap_4
XFILLER_76_797 VPWR VGND sg13g2_decap_8
XFILLER_64_959 VPWR VGND sg13g2_fill_1
XFILLER_48_499 VPWR VGND sg13g2_decap_4
XFILLER_35_105 VPWR VGND sg13g2_decap_8
X_14854_ _00655_ VGND VPWR _01378_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[5\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_1
XFILLER_17_831 VPWR VGND sg13g2_decap_8
X_14785_ _00586_ VGND VPWR _01309_ acc_sub.y\[14\] clknet_leaf_40_clk sg13g2_dfrbpq_1
XFILLER_91_778 VPWR VGND sg13g2_fill_1
X_13805_ VPWR _00356_ net73 VGND sg13g2_inv_1
XFILLER_63_458 VPWR VGND sg13g2_decap_8
X_11997_ _05851_ _05828_ _05826_ VPWR VGND sg13g2_xnor2_1
XFILLER_50_119 VPWR VGND sg13g2_decap_8
XFILLER_45_91 VPWR VGND sg13g2_decap_8
XFILLER_44_661 VPWR VGND sg13g2_decap_8
X_13736_ VPWR _00287_ net54 VGND sg13g2_inv_1
XFILLER_16_352 VPWR VGND sg13g2_decap_8
X_10948_ VGND VPWR _04743_ _04837_ _04954_ _04953_ sg13g2_a21oi_1
XFILLER_32_834 VPWR VGND sg13g2_decap_8
X_13667_ VPWR _00218_ net57 VGND sg13g2_inv_1
X_10879_ _04890_ _04889_ _04817_ VPWR VGND sg13g2_nand2_1
XFILLER_31_366 VPWR VGND sg13g2_decap_8
X_12618_ _06434_ _05339_ net1851 VPWR VGND sg13g2_nand2_1
X_13598_ VPWR _00149_ net62 VGND sg13g2_inv_1
X_12549_ _06363_ _06365_ _06366_ VPWR VGND sg13g2_nor2_1
XFILLER_8_573 VPWR VGND sg13g2_decap_8
X_14219_ VPWR _00770_ net105 VGND sg13g2_inv_1
XFILLER_6_63 VPWR VGND sg13g2_decap_8
XFILLER_125_482 VPWR VGND sg13g2_decap_8
XFILLER_113_600 VPWR VGND sg13g2_fill_1
XFILLER_113_655 VPWR VGND sg13g2_decap_4
XFILLER_98_366 VPWR VGND sg13g2_decap_8
XFILLER_4_790 VPWR VGND sg13g2_decap_8
XFILLER_112_176 VPWR VGND sg13g2_fill_2
X_09760_ _03647_ _03875_ _03876_ VPWR VGND sg13g2_nor2_1
XFILLER_86_517 VPWR VGND sg13g2_decap_8
X_09691_ _03805_ _03806_ _03807_ VPWR VGND sg13g2_nor2b_1
X_08711_ _02921_ VPWR _01334_ VGND net1814 _02920_ sg13g2_o21ai_1
XFILLER_20_0 VPWR VGND sg13g2_decap_8
XFILLER_94_550 VPWR VGND sg13g2_decap_8
X_08642_ _02862_ net1671 _02863_ VPWR VGND sg13g2_nor2_1
XFILLER_67_775 VPWR VGND sg13g2_decap_8
XFILLER_81_222 VPWR VGND sg13g2_decap_4
XFILLER_67_797 VPWR VGND sg13g2_fill_1
XFILLER_39_488 VPWR VGND sg13g2_fill_2
X_08573_ VPWR _02797_ acc_sum.op_sign_logic0.mantisa_b\[10\] VGND sg13g2_inv_1
XFILLER_82_756 VPWR VGND sg13g2_decap_4
XFILLER_54_458 VPWR VGND sg13g2_fill_2
XFILLER_63_981 VPWR VGND sg13g2_decap_8
XFILLER_41_119 VPWR VGND sg13g2_decap_8
XFILLER_23_801 VPWR VGND sg13g2_fill_1
XFILLER_23_812 VPWR VGND sg13g2_fill_2
XFILLER_23_823 VPWR VGND sg13g2_fill_1
XFILLER_25_28 VPWR VGND sg13g2_decap_8
X_07455_ VPWR _01778_ acc_sub.seg_reg0.q\[29\] VGND sg13g2_inv_1
XFILLER_50_686 VPWR VGND sg13g2_decap_8
X_07386_ _01732_ VPWR _01463_ VGND acc_sub.reg1en.d\[0\] _01731_ sg13g2_o21ai_1
XFILLER_109_928 VPWR VGND sg13g2_decap_8
X_09125_ VPWR _03305_ acc_sub.y\[8\] VGND sg13g2_inv_1
XFILLER_41_49 VPWR VGND sg13g2_decap_8
X_09056_ VGND VPWR net1786 _03241_ _03242_ _03136_ sg13g2_a21oi_1
XFILLER_108_427 VPWR VGND sg13g2_fill_1
X_08007_ net1843 _02273_ _02241_ _02274_ VPWR VGND sg13g2_nand3_1
XFILLER_104_622 VPWR VGND sg13g2_decap_4
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_104_666 VPWR VGND sg13g2_decap_8
XFILLER_104_633 VPWR VGND sg13g2_fill_1
X_08909_ _03014_ _03094_ _03096_ VPWR VGND sg13g2_nor2_2
XFILLER_106_75 VPWR VGND sg13g2_fill_1
XFILLER_66_35 VPWR VGND sg13g2_decap_8
XFILLER_57_230 VPWR VGND sg13g2_fill_1
X_09889_ fp16_res_pipe.op_sign_logic0.add_sub fp16_res_pipe.reg_add_sub.q\[0\] net1831
+ _01221_ VPWR VGND sg13g2_mux2_1
XFILLER_18_606 VPWR VGND sg13g2_decap_4
XFILLER_46_937 VPWR VGND sg13g2_fill_2
X_11920_ _05790_ VPWR _00994_ VGND net1881 _05789_ sg13g2_o21ai_1
XFILLER_122_63 VPWR VGND sg13g2_decap_8
X_11851_ VGND VPWR _05537_ _05664_ _05749_ _05663_ sg13g2_a21oi_1
X_14570_ _00371_ VGND VPWR net1846 fp16_sum_pipe.reg3en.q\[0\] clknet_leaf_97_clk
+ sg13g2_dfrbpq_2
X_10802_ _04814_ _03576_ _04780_ VPWR VGND sg13g2_xnor2_1
X_11782_ _05685_ _05684_ _05613_ _05490_ _05444_ VPWR VGND sg13g2_a22oi_1
XFILLER_14_812 VPWR VGND sg13g2_decap_4
XFILLER_26_683 VPWR VGND sg13g2_fill_2
X_13521_ VPWR _00072_ net83 VGND sg13g2_inv_1
XFILLER_13_333 VPWR VGND sg13g2_fill_1
XFILLER_14_867 VPWR VGND sg13g2_decap_8
X_10733_ net1824 fp16_res_pipe.add_renorm0.mantisa\[10\] _04746_ VPWR VGND sg13g2_nor2_2
XFILLER_25_182 VPWR VGND sg13g2_decap_8
XFILLER_41_653 VPWR VGND sg13g2_decap_8
XFILLER_51_1011 VPWR VGND sg13g2_fill_2
X_13452_ _07105_ VPWR _00778_ VGND _06925_ net1754 sg13g2_o21ai_1
X_10664_ _04677_ net1710 _04675_ VPWR VGND sg13g2_nand2_1
X_12403_ _06249_ _06248_ _06181_ VPWR VGND sg13g2_nand2_1
X_13383_ _07068_ net1695 sipo.word\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_40_196 VPWR VGND sg13g2_decap_4
X_10595_ _04610_ VPWR _01139_ VGND net1933 _02269_ sg13g2_o21ai_1
XFILLER_127_736 VPWR VGND sg13g2_decap_8
XFILLER_126_224 VPWR VGND sg13g2_decap_8
X_12334_ VPWR _06180_ _06179_ VGND sg13g2_inv_1
XFILLER_108_972 VPWR VGND sg13g2_decap_8
X_14004_ VPWR _00555_ net77 VGND sg13g2_inv_1
X_12265_ VPWR _06111_ _06110_ VGND sg13g2_inv_1
XFILLER_5_587 VPWR VGND sg13g2_decap_4
XFILLER_123_953 VPWR VGND sg13g2_decap_8
XFILLER_122_430 VPWR VGND sg13g2_decap_8
XFILLER_107_493 VPWR VGND sg13g2_decap_8
X_12196_ _06039_ fpmul.reg_b_out\[4\] _06037_ _06042_ VPWR VGND sg13g2_nand3_1
XFILLER_122_463 VPWR VGND sg13g2_decap_8
X_11147_ _05117_ net1698 _05079_ VPWR VGND sg13g2_nand2_1
XFILLER_68_539 VPWR VGND sg13g2_fill_2
XFILLER_68_528 VPWR VGND sg13g2_decap_8
XFILLER_96_859 VPWR VGND sg13g2_decap_8
XFILLER_95_369 VPWR VGND sg13g2_fill_1
X_11078_ _05055_ acc_sum.exp_mant_logic0.a\[12\] _05052_ _04993_ acc_sum.seg_reg0.q\[27\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_0_292 VPWR VGND sg13g2_decap_8
X_14906_ _00707_ VGND VPWR _01426_ acc_sub.op_sign_logic0.mantisa_a\[5\] clknet_leaf_68_clk
+ sg13g2_dfrbpq_2
XFILLER_37_959 VPWR VGND sg13g2_decap_8
XFILLER_36_436 VPWR VGND sg13g2_fill_2
X_10029_ _04116_ _04051_ _04117_ VPWR VGND sg13g2_nor2_1
X_14837_ _00638_ VGND VPWR _01361_ state\[3\] clknet_leaf_52_clk sg13g2_dfrbpq_1
XFILLER_63_244 VPWR VGND sg13g2_decap_8
XFILLER_36_469 VPWR VGND sg13g2_fill_1
XFILLER_91_586 VPWR VGND sg13g2_decap_8
X_14768_ _00569_ VGND VPWR _01292_ acc_sum.exp_mant_logic0.b\[13\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
XFILLER_51_439 VPWR VGND sg13g2_decap_4
XFILLER_44_480 VPWR VGND sg13g2_decap_4
XFILLER_32_631 VPWR VGND sg13g2_decap_8
X_14699_ _00500_ VGND VPWR _01227_ acc_sum.y\[2\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_13719_ VPWR _00270_ net60 VGND sg13g2_inv_1
XFILLER_20_815 VPWR VGND sg13g2_fill_1
X_07240_ _01610_ VPWR _01611_ VGND _01517_ _01519_ sg13g2_o21ai_1
XFILLER_60_995 VPWR VGND sg13g2_decap_8
XFILLER_32_686 VPWR VGND sg13g2_decap_8
X_07171_ _01536_ _01542_ _01543_ VPWR VGND sg13g2_nor2_1
XFILLER_9_871 VPWR VGND sg13g2_decap_8
XFILLER_118_747 VPWR VGND sg13g2_decap_8
XFILLER_117_224 VPWR VGND sg13g2_decap_8
XFILLER_68_0 VPWR VGND sg13g2_decap_8
XFILLER_8_370 VPWR VGND sg13g2_decap_8
XFILLER_115_1005 VPWR VGND sg13g2_decap_8
XFILLER_114_986 VPWR VGND sg13g2_decap_8
X_09812_ VPWR _03925_ _03859_ VGND sg13g2_inv_1
XFILLER_101_614 VPWR VGND sg13g2_decap_8
XFILLER_87_837 VPWR VGND sg13g2_decap_4
XFILLER_86_336 VPWR VGND sg13g2_fill_1
XFILLER_86_325 VPWR VGND sg13g2_decap_8
X_09743_ _03859_ _03855_ _03858_ VPWR VGND sg13g2_nand2_1
X_09674_ _03790_ _03789_ acc_sum.add_renorm0.exp\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_28_959 VPWR VGND sg13g2_decap_8
X_08625_ VPWR _02847_ _02846_ VGND sg13g2_inv_1
XFILLER_82_542 VPWR VGND sg13g2_decap_8
XFILLER_55_756 VPWR VGND sg13g2_decap_8
XFILLER_43_907 VPWR VGND sg13g2_decap_8
XFILLER_36_49 VPWR VGND sg13g2_decap_8
X_08556_ _02777_ _02779_ _02780_ VPWR VGND sg13g2_nor2_1
XFILLER_82_597 VPWR VGND sg13g2_decap_8
XFILLER_70_715 VPWR VGND sg13g2_decap_8
XFILLER_55_789 VPWR VGND sg13g2_decap_8
X_07507_ _01829_ _01828_ _01807_ VPWR VGND sg13g2_nand2b_1
XFILLER_23_620 VPWR VGND sg13g2_decap_8
X_08487_ _02663_ _02661_ _02715_ VPWR VGND sg13g2_nor2_1
XFILLER_51_962 VPWR VGND sg13g2_decap_8
X_07438_ fpdiv.divider0.divisor_reg\[7\] net1749 _01769_ VPWR VGND sg13g2_nor2_1
XFILLER_11_826 VPWR VGND sg13g2_fill_2
XFILLER_22_163 VPWR VGND sg13g2_decap_4
X_07369_ _01722_ net1799 acc_sub.seg_reg0.q\[23\] VPWR VGND sg13g2_nand2_1
XFILLER_6_307 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_fill_1
X_09108_ net1787 _03287_ _03285_ _03290_ VPWR VGND _03289_ sg13g2_nand4_1
XFILLER_108_246 VPWR VGND sg13g2_decap_8
X_10380_ VGND VPWR _04428_ _04420_ _04430_ _04427_ sg13g2_a21oi_1
XFILLER_124_739 VPWR VGND sg13g2_decap_8
X_09039_ _03225_ net1790 acc_sub.add_renorm0.exp\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_123_238 VPWR VGND sg13g2_decap_8
XFILLER_117_63 VPWR VGND sg13g2_decap_8
XFILLER_89_130 VPWR VGND sg13g2_fill_1
X_12050_ VPWR _05896_ _05895_ VGND sg13g2_inv_1
XFILLER_2_535 VPWR VGND sg13g2_decap_8
XFILLER_105_986 VPWR VGND sg13g2_decap_8
XFILLER_77_303 VPWR VGND sg13g2_fill_2
XFILLER_77_45 VPWR VGND sg13g2_decap_8
X_11001_ _04986_ VPWR _01109_ VGND net1929 _02459_ sg13g2_o21ai_1
XFILLER_77_347 VPWR VGND sg13g2_decap_8
XFILLER_77_67 VPWR VGND sg13g2_decap_8
XFILLER_77_56 VPWR VGND sg13g2_fill_1
XFILLER_120_967 VPWR VGND sg13g2_decap_8
XFILLER_93_807 VPWR VGND sg13g2_decap_8
XFILLER_86_870 VPWR VGND sg13g2_fill_2
XFILLER_58_550 VPWR VGND sg13g2_fill_1
XFILLER_46_701 VPWR VGND sg13g2_decap_8
XFILLER_19_915 VPWR VGND sg13g2_decap_8
X_12952_ _06724_ _06723_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_45_211 VPWR VGND sg13g2_decap_8
XFILLER_100_691 VPWR VGND sg13g2_decap_8
X_11903_ fpmul.seg_reg0.q\[47\] fpmul.reg_a_out\[8\] net1876 _01001_ VPWR VGND sg13g2_mux2_1
XFILLER_93_99 VPWR VGND sg13g2_fill_1
X_12883_ _00013_ net1731 net1702 _06660_ VPWR VGND sg13g2_nand3_1
XFILLER_60_203 VPWR VGND sg13g2_fill_1
X_14622_ _00423_ VGND VPWR _01154_ fp16_sum_pipe.add_renorm0.exp\[1\] clknet_leaf_111_clk
+ sg13g2_dfrbpq_2
XFILLER_27_981 VPWR VGND sg13g2_decap_8
XFILLER_33_428 VPWR VGND sg13g2_decap_8
X_11834_ _05444_ _05598_ _05733_ VPWR VGND sg13g2_nor2_1
X_14553_ _00354_ VGND VPWR _01089_ acc_sum.op_sign_logic0.mantisa_a\[5\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_11765_ _05656_ _05659_ _05668_ _05669_ VPWR VGND sg13g2_nor3_1
X_13504_ VPWR _00055_ net88 VGND sg13g2_inv_1
X_14484_ _00285_ VGND VPWR _01022_ add_result\[9\] clknet_leaf_99_clk sg13g2_dfrbpq_2
XFILLER_41_472 VPWR VGND sg13g2_fill_1
XFILLER_9_112 VPWR VGND sg13g2_decap_8
X_10716_ _04729_ _04675_ _04666_ _04670_ _04647_ VPWR VGND sg13g2_a22oi_1
X_13435_ _07096_ VPWR _00786_ VGND _06941_ net1720 sg13g2_o21ai_1
XFILLER_42_70 VPWR VGND sg13g2_decap_8
X_10647_ _04654_ _04658_ _04660_ VPWR VGND sg13g2_nor2_1
XFILLER_10_870 VPWR VGND sg13g2_decap_8
XFILLER_127_555 VPWR VGND sg13g2_decap_8
X_13366_ _07059_ net1696 sipo.word\[15\] VPWR VGND sg13g2_nand2_1
XFILLER_61_7 VPWR VGND sg13g2_fill_2
X_10578_ _04602_ acc_sub.x2\[10\] net1931 VPWR VGND sg13g2_nand2_1
XFILLER_115_739 VPWR VGND sg13g2_decap_8
X_13297_ _07010_ sipo.word\[3\] VPWR VGND sg13g2_inv_2
X_12317_ _06163_ net1857 net1868 VPWR VGND sg13g2_nand2_1
XFILLER_6_885 VPWR VGND sg13g2_decap_8
XFILLER_114_249 VPWR VGND sg13g2_decap_8
X_12248_ _06094_ net1869 _06093_ VPWR VGND sg13g2_xnor2_1
XFILLER_47_5 VPWR VGND sg13g2_decap_8
XFILLER_123_750 VPWR VGND sg13g2_decap_8
XFILLER_111_901 VPWR VGND sg13g2_decap_8
XFILLER_69_815 VPWR VGND sg13g2_decap_8
XFILLER_110_433 VPWR VGND sg13g2_decap_8
XFILLER_95_111 VPWR VGND sg13g2_fill_2
X_12179_ _06025_ fpmul.reg_b_out\[4\] VPWR VGND sg13g2_inv_2
XFILLER_3_42 VPWR VGND sg13g2_decap_8
XFILLER_111_978 VPWR VGND sg13g2_decap_8
XFILLER_110_466 VPWR VGND sg13g2_decap_4
XFILLER_95_133 VPWR VGND sg13g2_decap_8
XFILLER_95_199 VPWR VGND sg13g2_decap_8
XFILLER_36_211 VPWR VGND sg13g2_fill_2
X_08410_ VPWR _02645_ fpdiv.divider0.counter\[2\] VGND sg13g2_inv_1
XFILLER_92_873 VPWR VGND sg13g2_decap_4
XFILLER_91_361 VPWR VGND sg13g2_decap_8
XFILLER_52_715 VPWR VGND sg13g2_decap_8
XFILLER_51_203 VPWR VGND sg13g2_decap_8
XFILLER_36_277 VPWR VGND sg13g2_decap_8
X_09390_ VGND VPWR _03536_ _03397_ _03537_ _03518_ sg13g2_a21oi_1
X_08341_ sipo.word\[6\] sipo.word\[5\] sipo.word\[7\] _02586_ VPWR VGND sipo.word\[4\]
+ sg13g2_nand4_1
XFILLER_60_770 VPWR VGND sg13g2_fill_1
XFILLER_33_995 VPWR VGND sg13g2_decap_8
X_08272_ _02518_ _02520_ _02521_ VPWR VGND sg13g2_nor2_1
XFILLER_20_601 VPWR VGND sg13g2_decap_8
XFILLER_32_461 VPWR VGND sg13g2_fill_2
X_07223_ VGND VPWR _01591_ _01594_ _01595_ _01492_ sg13g2_a21oi_1
X_07154_ acc_sub.op_sign_logic0.mantisa_a\[6\] _01525_ _01526_ VPWR VGND sg13g2_nor2_2
XFILLER_118_588 VPWR VGND sg13g2_decap_8
XFILLER_102_923 VPWR VGND sg13g2_decap_8
Xfanout102 net104 net102 VPWR VGND sg13g2_buf_1
Xfanout113 net128 net113 VPWR VGND sg13g2_buf_1
Xfanout135 net136 net135 VPWR VGND sg13g2_buf_1
XFILLER_114_783 VPWR VGND sg13g2_decap_8
XFILLER_101_433 VPWR VGND sg13g2_decap_8
XFILLER_101_400 VPWR VGND sg13g2_decap_4
XFILLER_99_483 VPWR VGND sg13g2_fill_2
Xfanout124 net127 net124 VPWR VGND sg13g2_buf_2
XFILLER_59_314 VPWR VGND sg13g2_decap_8
XFILLER_87_689 VPWR VGND sg13g2_decap_8
XFILLER_59_369 VPWR VGND sg13g2_fill_2
XFILLER_59_358 VPWR VGND sg13g2_decap_4
XFILLER_47_26 VPWR VGND sg13g2_decap_8
X_07987_ _02256_ VPWR _01386_ VGND _02210_ _02248_ sg13g2_o21ai_1
X_09726_ _03842_ _03677_ _03680_ VPWR VGND sg13g2_nand2_1
XFILLER_28_712 VPWR VGND sg13g2_decap_8
XFILLER_103_32 VPWR VGND sg13g2_decap_8
X_09657_ _03773_ _03740_ _03774_ VPWR VGND sg13g2_and2_1
XFILLER_43_704 VPWR VGND sg13g2_decap_8
XFILLER_27_255 VPWR VGND sg13g2_decap_8
X_09588_ _03705_ net1805 acc_sum.add_renorm0.mantisa\[6\] VPWR VGND sg13g2_nand2_1
X_08608_ _02830_ VPWR _02831_ VGND _02780_ _02829_ sg13g2_o21ai_1
XFILLER_63_58 VPWR VGND sg13g2_decap_8
X_08539_ VPWR _02763_ acc_sum.op_sign_logic0.mantisa_a\[1\] VGND sg13g2_inv_1
XFILLER_23_450 VPWR VGND sg13g2_decap_8
XFILLER_51_770 VPWR VGND sg13g2_decap_8
X_11550_ _05454_ VPWR _05455_ VGND _05451_ _05439_ sg13g2_o21ai_1
XFILLER_24_995 VPWR VGND sg13g2_decap_8
XFILLER_10_133 VPWR VGND sg13g2_decap_8
X_10501_ _04545_ net1670 _04538_ VPWR VGND sg13g2_nand2_1
X_11481_ VPWR _05393_ fpdiv.divider0.divisor\[10\] VGND sg13g2_inv_1
X_13220_ _06947_ VPWR _00852_ VGND _06897_ _06880_ sg13g2_o21ai_1
XFILLER_6_126 VPWR VGND sg13g2_decap_8
XFILLER_11_689 VPWR VGND sg13g2_decap_8
X_10432_ VGND VPWR _04477_ _04478_ _04481_ _04480_ sg13g2_a21oi_1
XFILLER_88_11 VPWR VGND sg13g2_fill_2
X_13151_ VPWR _06897_ sipo.bit_counter\[2\] VGND sg13g2_inv_1
X_10363_ VPWR _04413_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[0\] VGND sg13g2_inv_1
XFILLER_12_84 VPWR VGND sg13g2_decap_8
XFILLER_124_536 VPWR VGND sg13g2_fill_2
X_13082_ _06846_ VPWR _00889_ VGND net1861 _06621_ sg13g2_o21ai_1
X_12102_ _05948_ _05892_ _05895_ VPWR VGND sg13g2_nand2_1
XFILLER_3_833 VPWR VGND sg13g2_decap_8
XFILLER_2_310 VPWR VGND sg13g2_fill_1
XFILLER_88_77 VPWR VGND sg13g2_decap_8
XFILLER_88_66 VPWR VGND sg13g2_fill_2
XFILLER_78_601 VPWR VGND sg13g2_fill_1
X_12033_ _00970_ _05878_ _05879_ _05877_ _05876_ VPWR VGND sg13g2_a22oi_1
X_10294_ _04329_ _04227_ _04362_ VPWR VGND sg13g2_nor2_1
XFILLER_120_764 VPWR VGND sg13g2_decap_8
XFILLER_66_829 VPWR VGND sg13g2_decap_8
XFILLER_66_818 VPWR VGND sg13g2_fill_1
XFILLER_92_114 VPWR VGND sg13g2_fill_2
XFILLER_92_103 VPWR VGND sg13g2_decap_8
XFILLER_65_339 VPWR VGND sg13g2_decap_8
XFILLER_65_317 VPWR VGND sg13g2_decap_8
XFILLER_59_870 VPWR VGND sg13g2_decap_8
XFILLER_58_380 VPWR VGND sg13g2_fill_1
X_13984_ VPWR _00535_ net25 VGND sg13g2_inv_1
X_12935_ _06707_ _06706_ fp16_sum_pipe.reg1en.d\[0\] _06708_ VPWR VGND sg13g2_a21o_2
XFILLER_46_586 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_18_266 VPWR VGND sg13g2_decap_8
X_12866_ _06645_ _06644_ fpmul.reg1en.d\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_18_288 VPWR VGND sg13g2_decap_8
XFILLER_61_556 VPWR VGND sg13g2_decap_8
X_11817_ _01024_ _05716_ _05717_ VPWR VGND sg13g2_nand2_1
XFILLER_15_973 VPWR VGND sg13g2_decap_8
X_14605_ _00406_ VGND VPWR _01137_ fp16_sum_pipe.exp_mant_logic0.a\[0\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_2
X_14536_ _00337_ VGND VPWR _01072_ fpdiv.div_out\[11\] clknet_leaf_77_clk sg13g2_dfrbpq_2
X_12797_ VGND VPWR net1935 add_result\[14\] _06581_ net1943 sg13g2_a21oi_1
XFILLER_14_472 VPWR VGND sg13g2_decap_8
XFILLER_119_308 VPWR VGND sg13g2_fill_1
X_11748_ VGND VPWR _05581_ net1839 _05652_ _05651_ sg13g2_a21oi_1
X_14467_ _00268_ VGND VPWR _01006_ fpmul.seg_reg0.q\[52\] clknet_leaf_125_clk sg13g2_dfrbpq_1
X_11679_ _05441_ _05440_ _05583_ VPWR VGND sg13g2_nor2_2
XFILLER_30_976 VPWR VGND sg13g2_decap_8
X_14398_ _00199_ VGND VPWR _00937_ div_result\[11\] clknet_leaf_89_clk sg13g2_dfrbpq_1
X_13418_ _07088_ net1722 instr\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_127_385 VPWR VGND sg13g2_decap_8
XFILLER_115_525 VPWR VGND sg13g2_fill_2
XFILLER_115_514 VPWR VGND sg13g2_decap_8
Xplace1805 acc_sum.add_renorm0.mantisa\[11\] net1805 VPWR VGND sg13g2_buf_2
Xplace1816 acc_sum.reg2en.q\[0\] net1816 VPWR VGND sg13g2_buf_2
X_13349_ _07048_ VPWR _00824_ VGND _06999_ net1723 sg13g2_o21ai_1
Xplace1827 fp16_res_pipe.exp_mant_logic0.a\[6\] net1827 VPWR VGND sg13g2_buf_2
Xplace1849 net1848 net1849 VPWR VGND sg13g2_buf_2
Xplace1838 fp16_sum_pipe.add_renorm0.mantisa\[11\] net1838 VPWR VGND sg13g2_buf_2
XFILLER_102_208 VPWR VGND sg13g2_decap_8
XFILLER_97_921 VPWR VGND sg13g2_decap_8
X_08890_ _03076_ _03057_ _03077_ VPWR VGND sg13g2_nor2b_1
XFILLER_68_111 VPWR VGND sg13g2_decap_8
X_07910_ VPWR _02185_ _02184_ VGND sg13g2_inv_1
X_07841_ _02137_ _02136_ net1640 VPWR VGND sg13g2_nand2_1
XFILLER_96_453 VPWR VGND sg13g2_decap_8
XFILLER_68_133 VPWR VGND sg13g2_decap_8
XFILLER_29_509 VPWR VGND sg13g2_decap_8
XFILLER_111_775 VPWR VGND sg13g2_decap_8
XFILLER_97_998 VPWR VGND sg13g2_decap_8
X_07772_ _02073_ acc_sub.exp_mant_logic0.b\[4\] VPWR VGND sg13g2_inv_2
XFILLER_83_103 VPWR VGND sg13g2_decap_8
XFILLER_56_317 VPWR VGND sg13g2_decap_8
X_09511_ acc_sum.add_renorm0.mantisa\[10\] _03627_ _03628_ VPWR VGND sg13g2_nor2_2
XFILLER_83_147 VPWR VGND sg13g2_fill_1
XFILLER_37_531 VPWR VGND sg13g2_fill_2
XFILLER_65_862 VPWR VGND sg13g2_decap_4
XFILLER_37_564 VPWR VGND sg13g2_decap_4
XFILLER_25_726 VPWR VGND sg13g2_decap_8
XFILLER_80_843 VPWR VGND sg13g2_fill_1
X_09442_ _03580_ fp16_res_pipe.add_renorm0.exp\[4\] VPWR VGND sg13g2_inv_2
X_09373_ _03389_ _03494_ _03522_ VPWR VGND sg13g2_nor2_1
X_08324_ _02568_ _02562_ _02569_ VPWR VGND sg13g2_nor2_1
XFILLER_40_729 VPWR VGND sg13g2_fill_1
XFILLER_33_770 VPWR VGND sg13g2_fill_2
XFILLER_21_910 VPWR VGND sg13g2_decap_8
XFILLER_33_28 VPWR VGND sg13g2_decap_8
XFILLER_20_420 VPWR VGND sg13g2_fill_2
X_08255_ _01367_ _02504_ _02505_ VPWR VGND sg13g2_nand2_1
XFILLER_20_475 VPWR VGND sg13g2_decap_8
XFILLER_21_987 VPWR VGND sg13g2_decap_8
XFILLER_119_842 VPWR VGND sg13g2_decap_8
X_07206_ VPWR _01578_ _01577_ VGND sg13g2_inv_1
X_08186_ _02444_ net1774 fp16_sum_pipe.op_sign_logic0.mantisa_a\[1\] VPWR VGND sg13g2_nand2_1
X_07137_ VPWR _01509_ acc_sub.op_sign_logic0.mantisa_a\[9\] VGND sg13g2_inv_1
XFILLER_109_7 VPWR VGND sg13g2_decap_8
XFILLER_0_814 VPWR VGND sg13g2_decap_8
XFILLER_58_14 VPWR VGND sg13g2_decap_8
XFILLER_102_742 VPWR VGND sg13g2_decap_8
XFILLER_101_230 VPWR VGND sg13g2_decap_4
XFILLER_75_604 VPWR VGND sg13g2_decap_8
XFILLER_114_42 VPWR VGND sg13g2_decap_8
XFILLER_102_786 VPWR VGND sg13g2_decap_4
XFILLER_47_306 VPWR VGND sg13g2_decap_4
XFILLER_28_531 VPWR VGND sg13g2_fill_2
X_09709_ net1769 VPWR _03825_ VGND _03795_ _03823_ sg13g2_o21ai_1
X_10981_ _04976_ VPWR _01119_ VGND net1926 _02463_ sg13g2_o21ai_1
XFILLER_83_681 VPWR VGND sg13g2_decap_8
X_12720_ _06526_ _06525_ _06513_ VPWR VGND sg13g2_nand2_1
XFILLER_15_203 VPWR VGND sg13g2_decap_4
XFILLER_16_759 VPWR VGND sg13g2_decap_8
XFILLER_82_191 VPWR VGND sg13g2_decap_8
X_12651_ _06416_ _06466_ _06467_ VPWR VGND sg13g2_nor2_1
XFILLER_71_876 VPWR VGND sg13g2_fill_2
XFILLER_43_567 VPWR VGND sg13g2_decap_8
XFILLER_15_236 VPWR VGND sg13g2_fill_2
XFILLER_15_269 VPWR VGND sg13g2_fill_1
XFILLER_70_397 VPWR VGND sg13g2_fill_1
XFILLER_12_932 VPWR VGND sg13g2_decap_8
X_11602_ _05482_ _05468_ _05507_ VPWR VGND sg13g2_nor2_1
X_12582_ _06377_ VPWR _06398_ VGND _05370_ fpdiv.reg_b_out\[7\] sg13g2_o21ai_1
XFILLER_11_442 VPWR VGND sg13g2_fill_1
XFILLER_90_89 VPWR VGND sg13g2_decap_8
X_14321_ _00122_ VGND VPWR _00864_ sipo.word\[9\] clknet_leaf_14_clk sg13g2_dfrbpq_2
XFILLER_7_402 VPWR VGND sg13g2_fill_2
X_11533_ _05436_ _05398_ _05419_ _05437_ _05438_ VPWR VGND sg13g2_nor4_1
XFILLER_99_21 VPWR VGND sg13g2_fill_2
X_14252_ _00053_ VGND VPWR _00803_ acc_sub.x2\[1\] clknet_leaf_50_clk sg13g2_dfrbpq_2
X_11464_ fpdiv.reg_b_out\[15\] fp16_res_pipe.x2\[15\] net1942 _01044_ VPWR VGND sg13g2_mux2_1
XFILLER_8_958 VPWR VGND sg13g2_decap_8
XFILLER_125_823 VPWR VGND sg13g2_decap_8
XFILLER_109_374 VPWR VGND sg13g2_decap_4
XFILLER_99_54 VPWR VGND sg13g2_fill_1
X_13203_ _06936_ VPWR _00858_ VGND _06935_ net1714 sg13g2_o21ai_1
X_10415_ _04464_ VPWR _01173_ VGND net1846 _04389_ sg13g2_o21ai_1
XFILLER_124_322 VPWR VGND sg13g2_decap_8
XFILLER_99_87 VPWR VGND sg13g2_fill_1
X_14183_ VPWR _00734_ net131 VGND sg13g2_inv_1
X_11395_ _05341_ VPWR _01070_ VGND _05339_ fpdiv.divider0.en_r sg13g2_o21ai_1
XFILLER_3_630 VPWR VGND sg13g2_decap_4
X_13134_ VPWR _06886_ _06885_ VGND sg13g2_inv_1
XFILLER_2_140 VPWR VGND sg13g2_decap_8
X_10346_ VPWR _04396_ _04395_ VGND sg13g2_inv_1
XFILLER_124_388 VPWR VGND sg13g2_fill_2
XFILLER_97_239 VPWR VGND sg13g2_fill_2
X_13065_ _06829_ _06830_ _06831_ _06832_ _06833_ VPWR VGND sg13g2_nor4_1
XFILLER_3_696 VPWR VGND sg13g2_decap_4
XFILLER_3_674 VPWR VGND sg13g2_decap_8
X_10277_ _04347_ _04346_ net1636 VPWR VGND sg13g2_nand2_1
XFILLER_120_550 VPWR VGND sg13g2_fill_2
X_12016_ net1874 fpmul.seg_reg0.q\[20\] _05867_ VPWR VGND sg13g2_nor2_1
XFILLER_24_7 VPWR VGND sg13g2_decap_8
XFILLER_78_464 VPWR VGND sg13g2_fill_2
XFILLER_94_968 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_19_531 VPWR VGND sg13g2_decap_8
XFILLER_94_1003 VPWR VGND sg13g2_decap_8
XFILLER_93_489 VPWR VGND sg13g2_fill_2
XFILLER_93_467 VPWR VGND sg13g2_decap_8
XFILLER_47_873 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
X_13967_ VPWR _00518_ net7 VGND sg13g2_inv_1
XFILLER_80_139 VPWR VGND sg13g2_decap_8
X_12918_ _06691_ _06692_ _06682_ _00899_ VPWR VGND sg13g2_nand3_1
XFILLER_62_865 VPWR VGND sg13g2_decap_4
XFILLER_34_545 VPWR VGND sg13g2_fill_1
X_13898_ VPWR _00449_ net17 VGND sg13g2_inv_1
XFILLER_0_98 VPWR VGND sg13g2_decap_8
X_12849_ VGND VPWR acc\[10\] net1907 _06629_ fp16_res_pipe.reg1en.d\[0\] sg13g2_a21oi_1
XFILLER_9_63 VPWR VGND sg13g2_decap_8
XFILLER_119_105 VPWR VGND sg13g2_decap_8
X_14519_ _00320_ VGND VPWR _01055_ fpdiv.reg_a_out\[10\] clknet_leaf_54_clk sg13g2_dfrbpq_1
XFILLER_30_762 VPWR VGND sg13g2_decap_8
XFILLER_127_182 VPWR VGND sg13g2_decap_8
XFILLER_116_856 VPWR VGND sg13g2_decap_8
Xplace1635 _05151_ net1635 VPWR VGND sg13g2_buf_2
XFILLER_50_0 VPWR VGND sg13g2_decap_8
Xplace1646 _01949_ net1646 VPWR VGND sg13g2_buf_2
Xplace1668 _02865_ net1668 VPWR VGND sg13g2_buf_2
XFILLER_89_707 VPWR VGND sg13g2_fill_2
Xplace1657 _02378_ net1657 VPWR VGND sg13g2_buf_2
X_09991_ _04079_ _04011_ _04014_ VPWR VGND sg13g2_nand2_1
X_08942_ _03127_ _03128_ _03126_ _03129_ VPWR VGND sg13g2_nand3_1
XFILLER_103_528 VPWR VGND sg13g2_decap_8
Xplace1679 _06962_ net1679 VPWR VGND sg13g2_buf_2
XFILLER_69_453 VPWR VGND sg13g2_decap_8
X_08873_ _03027_ _03031_ _03060_ VPWR VGND sg13g2_nor2_1
XFILLER_97_795 VPWR VGND sg13g2_decap_8
XFILLER_96_272 VPWR VGND sg13g2_fill_1
XFILLER_69_475 VPWR VGND sg13g2_decap_4
XFILLER_56_103 VPWR VGND sg13g2_fill_1
XFILLER_28_28 VPWR VGND sg13g2_decap_8
X_07824_ _02121_ _02119_ _02120_ VPWR VGND sg13g2_nand2_1
XFILLER_85_957 VPWR VGND sg13g2_decap_8
XFILLER_69_497 VPWR VGND sg13g2_decap_8
XFILLER_56_147 VPWR VGND sg13g2_decap_4
XFILLER_71_106 VPWR VGND sg13g2_decap_8
XFILLER_44_309 VPWR VGND sg13g2_fill_1
XFILLER_38_862 VPWR VGND sg13g2_decap_8
X_07686_ _01995_ acc_sub.exp_mant_logic0.a\[4\] net1649 net1792 _01975_ VPWR VGND
+ sg13g2_a22oi_1
XFILLER_37_394 VPWR VGND sg13g2_decap_8
XFILLER_44_49 VPWR VGND sg13g2_decap_8
X_09425_ _03567_ VPWR _03568_ VGND _03410_ net1675 sg13g2_o21ai_1
XFILLER_53_898 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_25_589 VPWR VGND sg13g2_decap_8
XFILLER_100_33 VPWR VGND sg13g2_fill_1
X_09356_ VGND VPWR _03496_ _03436_ _03507_ _03435_ sg13g2_a21oi_1
X_09287_ VPWR _03441_ _03425_ VGND sg13g2_inv_1
X_08307_ _02552_ VPWR _02553_ VGND _02467_ _02427_ sg13g2_o21ai_1
XFILLER_21_751 VPWR VGND sg13g2_decap_4
XFILLER_21_773 VPWR VGND sg13g2_decap_8
X_08238_ _01369_ _02489_ _02490_ VPWR VGND sg13g2_nand2_1
XFILLER_5_906 VPWR VGND sg13g2_decap_8
XFILLER_125_119 VPWR VGND sg13g2_decap_8
XFILLER_119_650 VPWR VGND sg13g2_decap_8
XFILLER_107_801 VPWR VGND sg13g2_fill_2
XFILLER_118_182 VPWR VGND sg13g2_decap_8
XFILLER_109_42 VPWR VGND sg13g2_decap_8
XFILLER_4_427 VPWR VGND sg13g2_decap_8
X_10200_ _04276_ net1644 net1829 VPWR VGND sg13g2_nand2_1
X_08169_ _02260_ _02427_ _02428_ VPWR VGND sg13g2_nor2_1
XFILLER_107_889 VPWR VGND sg13g2_fill_1
XFILLER_69_46 VPWR VGND sg13g2_decap_8
X_11180_ _05143_ _05148_ _05138_ _05149_ VPWR VGND sg13g2_nand3_1
XFILLER_122_826 VPWR VGND sg13g2_decap_8
X_10131_ _04209_ _04212_ _04213_ VPWR VGND sg13g2_nor2_1
XFILLER_76_902 VPWR VGND sg13g2_decap_4
XFILLER_0_644 VPWR VGND sg13g2_decap_8
X_10062_ _04054_ _04149_ _04150_ VPWR VGND sg13g2_nor2_1
XFILLER_125_63 VPWR VGND sg13g2_decap_8
XFILLER_76_924 VPWR VGND sg13g2_fill_1
XFILLER_47_103 VPWR VGND sg13g2_decap_8
X_14870_ _00671_ VGND VPWR net1800 acc_sub.reg4en.q\[0\] clknet_leaf_45_clk sg13g2_dfrbpq_1
XFILLER_85_67 VPWR VGND sg13g2_decap_4
XFILLER_85_45 VPWR VGND sg13g2_fill_2
XFILLER_75_456 VPWR VGND sg13g2_decap_8
X_13821_ VPWR _00372_ net44 VGND sg13g2_inv_1
X_13752_ VPWR _00303_ net109 VGND sg13g2_inv_1
XFILLER_62_139 VPWR VGND sg13g2_fill_2
XFILLER_56_692 VPWR VGND sg13g2_decap_8
X_12703_ _06511_ _06453_ _06425_ VPWR VGND sg13g2_nand2_1
XFILLER_55_191 VPWR VGND sg13g2_fill_2
X_10964_ fp16_res_pipe.y\[6\] _04732_ net1835 _01127_ VPWR VGND sg13g2_mux2_1
X_13683_ VPWR _00234_ net62 VGND sg13g2_inv_1
XFILLER_31_504 VPWR VGND sg13g2_decap_8
XFILLER_31_515 VPWR VGND sg13g2_fill_2
X_10895_ _04737_ VPWR _04905_ VGND _04851_ _04904_ sg13g2_o21ai_1
X_12634_ VPWR _06450_ _06449_ VGND sg13g2_inv_1
XFILLER_70_194 VPWR VGND sg13g2_decap_8
XFILLER_86_9 VPWR VGND sg13g2_fill_1
X_12565_ _06381_ _06379_ _06380_ VPWR VGND sg13g2_xnor2_1
XFILLER_102_1007 VPWR VGND sg13g2_decap_8
X_14304_ _00105_ VGND VPWR _00848_ acc\[14\] clknet_leaf_49_clk sg13g2_dfrbpq_2
XFILLER_7_221 VPWR VGND sg13g2_fill_2
XFILLER_7_210 VPWR VGND sg13g2_decap_8
X_11516_ _05420_ VPWR _05421_ VGND net1841 _05419_ sg13g2_o21ai_1
X_12496_ _06331_ _06233_ _06239_ VPWR VGND sg13g2_xnor2_1
XFILLER_7_265 VPWR VGND sg13g2_fill_2
XFILLER_7_254 VPWR VGND sg13g2_decap_8
X_11447_ VPWR _05374_ fpdiv.divider0.dividend\[9\] VGND sg13g2_inv_1
X_14235_ _00036_ VGND VPWR _00786_ instr\[0\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_50_70 VPWR VGND sg13g2_decap_8
XFILLER_7_298 VPWR VGND sg13g2_decap_8
X_14166_ VPWR _00717_ net90 VGND sg13g2_inv_1
X_11378_ _05329_ _05328_ net1634 VPWR VGND sg13g2_nand2_1
XFILLER_4_972 VPWR VGND sg13g2_decap_8
XFILLER_113_837 VPWR VGND sg13g2_decap_8
X_13117_ _06783_ VPWR _06873_ VGND _06779_ _06868_ sg13g2_o21ai_1
X_10329_ _04382_ net1920 fp16_res_pipe.x2\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_124_196 VPWR VGND sg13g2_decap_8
XFILLER_112_358 VPWR VGND sg13g2_decap_8
XFILLER_79_740 VPWR VGND sg13g2_fill_2
X_14097_ VPWR _00648_ net41 VGND sg13g2_inv_1
XFILLER_94_721 VPWR VGND sg13g2_fill_1
XFILLER_78_261 VPWR VGND sg13g2_decap_8
XFILLER_78_250 VPWR VGND sg13g2_decap_4
X_13048_ _06748_ _06815_ _06816_ VPWR VGND sg13g2_nor2_1
XFILLER_66_423 VPWR VGND sg13g2_decap_8
XFILLER_82_905 VPWR VGND sg13g2_decap_8
XFILLER_67_979 VPWR VGND sg13g2_fill_2
X_07540_ _01858_ _01847_ acc_sub.exp_mant_logic0.a\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_47_670 VPWR VGND sg13g2_fill_2
XFILLER_90_960 VPWR VGND sg13g2_decap_8
XFILLER_35_843 VPWR VGND sg13g2_fill_2
XFILLER_34_342 VPWR VGND sg13g2_decap_4
X_07471_ acc_sub.exp_mant_logic0.b\[12\] _01729_ _01794_ VPWR VGND sg13g2_nor2_1
XFILLER_61_161 VPWR VGND sg13g2_decap_8
XFILLER_50_813 VPWR VGND sg13g2_fill_1
XFILLER_98_0 VPWR VGND sg13g2_decap_4
X_09210_ _03361_ _03364_ _03365_ VPWR VGND sg13g2_nor2_1
XFILLER_22_548 VPWR VGND sg13g2_decap_8
X_09141_ acc_sub.y\[7\] net1773 _03319_ _01302_ VPWR VGND sg13g2_a21o_1
X_09072_ VGND VPWR net1786 _03256_ _03257_ _03136_ sg13g2_a21oi_1
X_08023_ _02236_ VPWR _02289_ VGND _02200_ _02288_ sg13g2_o21ai_1
XFILLER_1_408 VPWR VGND sg13g2_decap_8
XFILLER_116_686 VPWR VGND sg13g2_decap_8
XFILLER_104_826 VPWR VGND sg13g2_decap_8
XFILLER_115_196 VPWR VGND sg13g2_decap_8
X_09974_ _04065_ _04052_ fp16_res_pipe.exp_mant_logic0.b\[8\] VPWR VGND sg13g2_nand2_1
X_08925_ acc_sub.seg_reg1.q\[21\] _03111_ _03112_ VPWR VGND sg13g2_nor2_1
XFILLER_85_721 VPWR VGND sg13g2_fill_2
XFILLER_39_49 VPWR VGND sg13g2_decap_8
XFILLER_97_592 VPWR VGND sg13g2_fill_1
XFILLER_58_957 VPWR VGND sg13g2_decap_8
X_07807_ VGND VPWR acc_sub.exp_mant_logic0.b\[3\] net1646 _02105_ _02104_ sg13g2_a21oi_1
XFILLER_72_404 VPWR VGND sg13g2_decap_8
XFILLER_57_478 VPWR VGND sg13g2_decap_8
X_08787_ VPWR _02974_ acc_sub.add_renorm0.mantisa\[9\] VGND sg13g2_inv_1
XFILLER_84_297 VPWR VGND sg13g2_fill_1
XFILLER_72_437 VPWR VGND sg13g2_decap_8
XFILLER_57_489 VPWR VGND sg13g2_fill_1
XFILLER_26_821 VPWR VGND sg13g2_decap_8
XFILLER_111_21 VPWR VGND sg13g2_decap_8
X_07738_ _02043_ _02006_ acc_sub.exp_mant_logic0.a\[4\] VPWR VGND sg13g2_nand2_1
XFILLER_37_180 VPWR VGND sg13g2_decap_4
X_07669_ _01979_ _01923_ VPWR VGND sg13g2_inv_2
XFILLER_81_971 VPWR VGND sg13g2_decap_8
XFILLER_40_301 VPWR VGND sg13g2_decap_4
XFILLER_26_898 VPWR VGND sg13g2_decap_8
XFILLER_111_98 VPWR VGND sg13g2_decap_4
XFILLER_80_492 VPWR VGND sg13g2_decap_8
XFILLER_71_47 VPWR VGND sg13g2_fill_1
XFILLER_71_36 VPWR VGND sg13g2_decap_8
XFILLER_52_194 VPWR VGND sg13g2_decap_4
X_10680_ _04664_ _04675_ _04692_ _04693_ VPWR VGND sg13g2_nand3_1
X_09408_ VGND VPWR _03552_ _03464_ _03553_ _03518_ sg13g2_a21oi_1
X_09339_ VGND VPWR _03490_ _03418_ _03491_ _03401_ sg13g2_a21oi_1
XFILLER_9_519 VPWR VGND sg13g2_decap_8
XFILLER_40_389 VPWR VGND sg13g2_fill_2
XFILLER_127_918 VPWR VGND sg13g2_decap_8
X_12350_ _06162_ VPWR _06196_ VGND _06065_ _06165_ sg13g2_o21ai_1
XFILLER_5_714 VPWR VGND sg13g2_decap_8
XFILLER_119_491 VPWR VGND sg13g2_fill_2
X_12281_ _06127_ _06124_ _06126_ VPWR VGND sg13g2_nand2_1
X_11301_ _01082_ _05258_ _05259_ VPWR VGND sg13g2_nand2_1
XFILLER_5_747 VPWR VGND sg13g2_decap_4
XFILLER_4_224 VPWR VGND sg13g2_decap_8
X_14020_ VPWR _00571_ net87 VGND sg13g2_inv_1
X_11232_ _05190_ _05195_ _05196_ _05197_ VPWR VGND sg13g2_nor3_1
XFILLER_4_257 VPWR VGND sg13g2_decap_8
XFILLER_4_246 VPWR VGND sg13g2_fill_2
XFILLER_106_174 VPWR VGND sg13g2_fill_1
X_11163_ _05024_ _05131_ _05130_ _05132_ VPWR VGND sg13g2_nand3_1
XFILLER_1_920 VPWR VGND sg13g2_decap_8
XFILLER_121_133 VPWR VGND sg13g2_decap_8
X_10114_ _04196_ VPWR _04197_ VGND _03611_ _04156_ sg13g2_o21ai_1
XFILLER_110_829 VPWR VGND sg13g2_decap_8
XFILLER_96_77 VPWR VGND sg13g2_decap_8
XFILLER_95_507 VPWR VGND sg13g2_decap_8
X_11094_ _05065_ _05066_ _05064_ _01096_ VPWR VGND sg13g2_nand3_1
XFILLER_49_924 VPWR VGND sg13g2_decap_8
XFILLER_0_463 VPWR VGND sg13g2_decap_8
XFILLER_1_997 VPWR VGND sg13g2_decap_8
X_14922_ _00723_ VGND VPWR _01442_ acc_sub.op_sign_logic0.s_a clknet_leaf_42_clk sg13g2_dfrbpq_1
XFILLER_103_892 VPWR VGND sg13g2_fill_1
XFILLER_75_220 VPWR VGND sg13g2_decap_8
X_10045_ net1703 VPWR _04133_ VGND _04130_ _04131_ sg13g2_o21ai_1
XFILLER_64_927 VPWR VGND sg13g2_decap_8
X_14853_ _00654_ VGND VPWR _01377_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[4\] clknet_leaf_114_clk
+ sg13g2_dfrbpq_2
X_13804_ VPWR _00355_ net73 VGND sg13g2_inv_1
XFILLER_75_275 VPWR VGND sg13g2_fill_1
XFILLER_64_938 VPWR VGND sg13g2_fill_2
XFILLER_63_437 VPWR VGND sg13g2_decap_4
XFILLER_57_990 VPWR VGND sg13g2_fill_2
X_14784_ _00585_ VGND VPWR _01308_ acc_sub.y\[13\] clknet_leaf_37_clk sg13g2_dfrbpq_1
X_11996_ _05849_ VPWR _05850_ VGND _05830_ _05831_ sg13g2_o21ai_1
XFILLER_16_331 VPWR VGND sg13g2_decap_4
XFILLER_17_843 VPWR VGND sg13g2_decap_4
X_13735_ VPWR _00286_ net68 VGND sg13g2_inv_1
XFILLER_45_70 VPWR VGND sg13g2_decap_8
XFILLER_17_898 VPWR VGND sg13g2_decap_8
X_10947_ fp16_res_pipe.seg_reg1.q\[21\] VPWR _04953_ VGND _04837_ _04774_ sg13g2_o21ai_1
XFILLER_31_301 VPWR VGND sg13g2_fill_1
X_13666_ VPWR _00217_ net57 VGND sg13g2_inv_1
XFILLER_43_183 VPWR VGND sg13g2_decap_4
XFILLER_31_334 VPWR VGND sg13g2_decap_8
X_12617_ _06428_ _06432_ _06433_ VPWR VGND sg13g2_nor2_1
X_10878_ _04889_ _04888_ _04797_ VPWR VGND sg13g2_nand2_1
Xclkbuf_4_14_0_clk clknet_0_clk clknet_4_14_0_clk VPWR VGND sg13g2_buf_8
X_13597_ VPWR _00148_ net110 VGND sg13g2_inv_1
XFILLER_118_929 VPWR VGND sg13g2_decap_8
X_12548_ _05387_ _05389_ _06364_ _06365_ VPWR VGND _05391_ sg13g2_nand4_1
XFILLER_117_439 VPWR VGND sg13g2_decap_8
X_12479_ VGND VPWR _06317_ net1872 _00963_ _06318_ sg13g2_a21oi_1
XFILLER_6_42 VPWR VGND sg13g2_decap_8
X_14218_ VPWR _00769_ net105 VGND sg13g2_inv_1
XFILLER_126_995 VPWR VGND sg13g2_decap_8
X_14149_ VPWR _00700_ net134 VGND sg13g2_inv_1
XFILLER_113_667 VPWR VGND sg13g2_decap_8
XFILLER_112_111 VPWR VGND sg13g2_decap_8
XFILLER_101_818 VPWR VGND sg13g2_decap_8
XFILLER_112_188 VPWR VGND sg13g2_fill_2
XFILLER_100_339 VPWR VGND sg13g2_fill_2
XFILLER_100_328 VPWR VGND sg13g2_decap_8
X_09690_ _03806_ acc_sum.add_renorm0.mantisa\[11\] acc_sum.add_renorm0.exp\[0\] VPWR
+ VGND sg13g2_nand2_1
X_08710_ _02921_ net1819 acc_sum.seg_reg0.q\[29\] VPWR VGND sg13g2_nand2_1
XFILLER_6_1013 VPWR VGND sg13g2_fill_1
XFILLER_94_562 VPWR VGND sg13g2_decap_4
X_08641_ VGND VPWR _02787_ _02790_ _02862_ _02733_ sg13g2_a21oi_1
XFILLER_67_754 VPWR VGND sg13g2_decap_8
XFILLER_66_231 VPWR VGND sg13g2_decap_8
XFILLER_55_927 VPWR VGND sg13g2_fill_1
XFILLER_55_916 VPWR VGND sg13g2_decap_8
XFILLER_13_0 VPWR VGND sg13g2_decap_8
XFILLER_55_949 VPWR VGND sg13g2_decap_8
X_08572_ acc_sum.op_sign_logic0.mantisa_b\[10\] _02795_ _02796_ VPWR VGND sg13g2_nor2_1
XFILLER_81_245 VPWR VGND sg13g2_decap_8
XFILLER_70_908 VPWR VGND sg13g2_fill_2
X_07523_ _01779_ _01843_ _01844_ VPWR VGND sg13g2_nor2_2
XFILLER_34_161 VPWR VGND sg13g2_decap_4
X_07454_ acc_sub.op_sign_logic0.add_sub acc_sub.reg_add_sub.q\[0\] acc_sub.reg1en.q\[0\]
+ _01440_ VPWR VGND sg13g2_mux2_1
XFILLER_62_481 VPWR VGND sg13g2_decap_4
XFILLER_109_907 VPWR VGND sg13g2_decap_8
X_07385_ _01732_ acc_sub.reg1en.d\[0\] acc\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_22_389 VPWR VGND sg13g2_fill_2
X_09124_ _03304_ VPWR _01304_ VGND net1801 _03294_ sg13g2_o21ai_1
X_09055_ _03241_ _03217_ _03240_ VPWR VGND sg13g2_xnor2_1
XFILLER_108_439 VPWR VGND sg13g2_decap_4
XFILLER_68_1008 VPWR VGND sg13g2_decap_4
X_08006_ _02272_ _02273_ VPWR VGND sg13g2_inv_4
XFILLER_117_984 VPWR VGND sg13g2_decap_8
XFILLER_89_323 VPWR VGND sg13g2_decap_8
XFILLER_104_645 VPWR VGND sg13g2_decap_8
XFILLER_103_122 VPWR VGND sg13g2_decap_8
XFILLER_106_54 VPWR VGND sg13g2_fill_2
XFILLER_106_43 VPWR VGND sg13g2_decap_8
XFILLER_89_378 VPWR VGND sg13g2_fill_1
XFILLER_77_518 VPWR VGND sg13g2_decap_8
X_09957_ net1766 _04051_ _04052_ VPWR VGND sg13g2_nor2_2
XFILLER_98_890 VPWR VGND sg13g2_fill_1
XFILLER_66_14 VPWR VGND sg13g2_decap_8
XFILLER_100_851 VPWR VGND sg13g2_fill_2
XFILLER_58_776 VPWR VGND sg13g2_fill_2
XFILLER_58_765 VPWR VGND sg13g2_fill_1
X_09888_ VGND VPWR net1831 _03985_ _01222_ _03986_ sg13g2_a21oi_1
X_08839_ _03026_ _03024_ _03025_ VPWR VGND sg13g2_nand2_1
XFILLER_85_595 VPWR VGND sg13g2_decap_8
XFILLER_57_275 VPWR VGND sg13g2_fill_2
XFILLER_122_42 VPWR VGND sg13g2_decap_8
XFILLER_73_779 VPWR VGND sg13g2_decap_8
XFILLER_73_757 VPWR VGND sg13g2_decap_4
XFILLER_57_297 VPWR VGND sg13g2_decap_8
X_11850_ net1837 _05746_ _05745_ _05748_ VPWR VGND _05747_ sg13g2_nand4_1
XFILLER_82_35 VPWR VGND sg13g2_decap_8
XFILLER_54_993 VPWR VGND sg13g2_fill_2
XFILLER_54_982 VPWR VGND sg13g2_decap_8
X_11781_ _05684_ _05611_ _05627_ VPWR VGND sg13g2_nand2_1
XFILLER_26_662 VPWR VGND sg13g2_decap_8
X_10801_ _04798_ _04812_ _04813_ VPWR VGND sg13g2_nor2_1
X_13520_ VPWR _00071_ net83 VGND sg13g2_inv_1
XFILLER_41_632 VPWR VGND sg13g2_decap_8
XFILLER_14_846 VPWR VGND sg13g2_decap_8
X_10732_ VGND VPWR _04739_ _04744_ _04745_ net1771 sg13g2_a21oi_1
XFILLER_25_161 VPWR VGND sg13g2_decap_8
XFILLER_9_316 VPWR VGND sg13g2_decap_8
XFILLER_13_356 VPWR VGND sg13g2_decap_8
X_13451_ _07105_ net1754 sipo.shift_reg\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_40_175 VPWR VGND sg13g2_decap_8
XFILLER_9_327 VPWR VGND sg13g2_fill_1
XFILLER_127_715 VPWR VGND sg13g2_decap_8
X_12402_ _06248_ _06183_ _06184_ VPWR VGND sg13g2_nand2_1
X_13382_ _07067_ VPWR _00810_ VGND _03601_ net1695 sg13g2_o21ai_1
X_10594_ _04610_ acc_sub.x2\[2\] net1934 VPWR VGND sg13g2_nand2_1
XFILLER_126_203 VPWR VGND sg13g2_decap_8
X_12333_ _06086_ _06178_ _06156_ _06179_ VPWR VGND sg13g2_nand3_1
XFILLER_108_951 VPWR VGND sg13g2_decap_8
XFILLER_123_932 VPWR VGND sg13g2_decap_8
X_14003_ VPWR _00554_ net79 VGND sg13g2_inv_1
Xoutput4 net4 miso VPWR VGND sg13g2_buf_1
X_12264_ VGND VPWR _06084_ _06108_ _06110_ _06109_ sg13g2_a21oi_1
XFILLER_122_442 VPWR VGND sg13g2_decap_4
X_11215_ net1663 _05180_ _05181_ VPWR VGND sg13g2_nor2b_2
X_12195_ _06041_ _06040_ _06025_ VPWR VGND sg13g2_nand2_1
XFILLER_96_838 VPWR VGND sg13g2_decap_8
X_11146_ _05115_ _05014_ _05116_ VPWR VGND sg13g2_xor2_1
XFILLER_68_507 VPWR VGND sg13g2_decap_8
XFILLER_89_890 VPWR VGND sg13g2_fill_1
XFILLER_49_732 VPWR VGND sg13g2_decap_8
XFILLER_0_271 VPWR VGND sg13g2_decap_8
XFILLER_0_260 VPWR VGND sg13g2_decap_8
X_14905_ _00706_ VGND VPWR _01425_ acc_sub.op_sign_logic0.mantisa_a\[4\] clknet_leaf_68_clk
+ sg13g2_dfrbpq_2
X_10028_ VGND VPWR _04081_ _04024_ _04116_ _04037_ sg13g2_a21oi_1
XFILLER_76_595 VPWR VGND sg13g2_fill_1
XFILLER_76_584 VPWR VGND sg13g2_fill_2
XFILLER_64_713 VPWR VGND sg13g2_decap_4
XFILLER_63_212 VPWR VGND sg13g2_fill_1
XFILLER_49_787 VPWR VGND sg13g2_decap_8
XFILLER_37_938 VPWR VGND sg13g2_decap_8
XFILLER_36_415 VPWR VGND sg13g2_decap_8
XFILLER_91_554 VPWR VGND sg13g2_decap_4
X_14836_ _00637_ VGND VPWR _01360_ state\[2\] clknet_leaf_51_clk sg13g2_dfrbpq_2
XFILLER_64_746 VPWR VGND sg13g2_decap_8
XFILLER_91_565 VPWR VGND sg13g2_decap_8
X_14767_ _00568_ VGND VPWR _01291_ acc_sum.exp_mant_logic0.b\[12\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
XFILLER_17_662 VPWR VGND sg13g2_fill_1
X_11979_ VPWR _05833_ _05832_ VGND sg13g2_inv_1
X_13718_ VPWR _00269_ net57 VGND sg13g2_inv_1
XFILLER_16_172 VPWR VGND sg13g2_decap_4
X_14698_ _00499_ VGND VPWR _01226_ acc_sum.y\[1\] clknet_leaf_47_clk sg13g2_dfrbpq_1
XFILLER_31_142 VPWR VGND sg13g2_decap_8
X_13649_ VPWR _00200_ net110 VGND sg13g2_inv_1
XFILLER_20_849 VPWR VGND sg13g2_fill_1
XFILLER_31_186 VPWR VGND sg13g2_decap_8
X_07170_ VPWR _01542_ _01541_ VGND sg13g2_inv_1
XFILLER_9_850 VPWR VGND sg13g2_decap_8
XFILLER_118_726 VPWR VGND sg13g2_decap_8
XFILLER_117_203 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_120_clk clknet_5_11__leaf_clk clknet_leaf_120_clk VPWR VGND sg13g2_buf_8
XFILLER_126_792 VPWR VGND sg13g2_decap_8
XFILLER_125_280 VPWR VGND sg13g2_decap_8
XFILLER_114_965 VPWR VGND sg13g2_decap_8
XFILLER_99_654 VPWR VGND sg13g2_decap_8
X_09811_ _03923_ VPWR _03924_ VGND _03647_ _03921_ sg13g2_o21ai_1
XFILLER_99_676 VPWR VGND sg13g2_fill_1
XFILLER_98_153 VPWR VGND sg13g2_fill_1
XFILLER_98_142 VPWR VGND sg13g2_decap_8
XFILLER_86_304 VPWR VGND sg13g2_decap_8
X_09742_ _03858_ _03857_ VPWR VGND sg13g2_inv_2
XFILLER_101_648 VPWR VGND sg13g2_fill_1
XFILLER_98_197 VPWR VGND sg13g2_decap_8
XFILLER_100_136 VPWR VGND sg13g2_decap_4
XFILLER_94_370 VPWR VGND sg13g2_decap_4
X_09673_ _02926_ _03788_ _03789_ VPWR VGND sg13g2_nor2_1
XFILLER_55_735 VPWR VGND sg13g2_decap_8
XFILLER_55_713 VPWR VGND sg13g2_fill_1
XFILLER_36_28 VPWR VGND sg13g2_decap_8
XFILLER_28_938 VPWR VGND sg13g2_decap_8
X_08624_ VGND VPWR _02845_ _02756_ _02846_ _02755_ sg13g2_a21oi_1
XFILLER_55_768 VPWR VGND sg13g2_decap_8
X_08555_ VPWR _02779_ _02778_ VGND sg13g2_inv_1
XFILLER_82_576 VPWR VGND sg13g2_fill_2
XFILLER_54_278 VPWR VGND sg13g2_fill_1
XFILLER_54_267 VPWR VGND sg13g2_fill_2
X_07506_ _01828_ _01827_ _01810_ VPWR VGND sg13g2_nand2_1
X_08486_ _02714_ VPWR _01352_ VGND net1705 _02713_ sg13g2_o21ai_1
XFILLER_22_142 VPWR VGND sg13g2_decap_8
X_07437_ VPWR _01768_ fpdiv.divider0.divisor\[7\] VGND sg13g2_inv_1
XFILLER_10_315 VPWR VGND sg13g2_decap_4
X_07368_ _01721_ acc_sub.add_renorm0.exp\[1\] VPWR VGND sg13g2_inv_2
XFILLER_22_186 VPWR VGND sg13g2_fill_1
X_09107_ _03097_ VPWR _03289_ VGND _03288_ _03208_ sg13g2_o21ai_1
XFILLER_108_214 VPWR VGND sg13g2_fill_2
X_07299_ _01664_ VPWR _01665_ VGND _01575_ net1667 sg13g2_o21ai_1
Xclkbuf_leaf_111_clk clknet_5_10__leaf_clk clknet_leaf_111_clk VPWR VGND sg13g2_buf_8
XFILLER_123_217 VPWR VGND sg13g2_decap_8
XFILLER_117_781 VPWR VGND sg13g2_decap_8
X_09038_ net1790 acc_sub.add_renorm0.exp\[0\] _03224_ VPWR VGND sg13g2_nor2_1
XFILLER_2_514 VPWR VGND sg13g2_decap_8
XFILLER_117_42 VPWR VGND sg13g2_decap_8
XFILLER_105_965 VPWR VGND sg13g2_decap_8
XFILLER_78_805 VPWR VGND sg13g2_decap_4
X_11000_ _04986_ fp16_res_pipe.x2\[4\] net1928 VPWR VGND sg13g2_nand2_1
XFILLER_120_946 VPWR VGND sg13g2_decap_8
XFILLER_92_329 VPWR VGND sg13g2_fill_2
X_12951_ _06722_ VPWR _06723_ VGND net1961 _06720_ sg13g2_o21ai_1
XFILLER_46_724 VPWR VGND sg13g2_fill_2
XFILLER_46_713 VPWR VGND sg13g2_fill_1
XFILLER_73_554 VPWR VGND sg13g2_decap_4
X_12882_ _06658_ _06659_ _06649_ _00902_ VPWR VGND sg13g2_nand3_1
X_11902_ fpmul.seg_reg0.q\[48\] fpmul.reg_a_out\[9\] net1876 _01002_ VPWR VGND sg13g2_mux2_1
XFILLER_18_448 VPWR VGND sg13g2_decap_4
XFILLER_93_78 VPWR VGND sg13g2_fill_2
XFILLER_73_587 VPWR VGND sg13g2_decap_8
XFILLER_34_919 VPWR VGND sg13g2_decap_8
XFILLER_27_960 VPWR VGND sg13g2_decap_8
X_14621_ _00422_ VGND VPWR _01153_ fp16_sum_pipe.add_renorm0.exp\[0\] clknet_leaf_111_clk
+ sg13g2_dfrbpq_2
X_11833_ _05732_ _05731_ _05720_ VPWR VGND sg13g2_nand2_1
XFILLER_33_407 VPWR VGND sg13g2_decap_4
XFILLER_54_790 VPWR VGND sg13g2_fill_2
XFILLER_14_632 VPWR VGND sg13g2_fill_1
X_14552_ _00353_ VGND VPWR _01088_ acc_sum.op_sign_logic0.mantisa_a\[4\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
XFILLER_60_259 VPWR VGND sg13g2_decap_8
X_11764_ VPWR _05668_ _05667_ VGND sg13g2_inv_1
X_13503_ VPWR _00054_ net89 VGND sg13g2_inv_1
X_14483_ _00284_ VGND VPWR _01021_ add_result\[8\] clknet_leaf_98_clk sg13g2_dfrbpq_2
X_10715_ _04658_ VPWR _04728_ VGND net1710 _04662_ sg13g2_o21ai_1
X_11695_ _05598_ _05444_ _05592_ _05599_ VPWR VGND sg13g2_nand3_1
X_13434_ _07096_ net1720 instr\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_127_534 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_102_clk clknet_5_15__leaf_clk clknet_leaf_102_clk VPWR VGND sg13g2_buf_8
X_10577_ _04601_ VPWR _01148_ VGND net1926 _02192_ sg13g2_o21ai_1
XFILLER_6_864 VPWR VGND sg13g2_decap_8
XFILLER_115_718 VPWR VGND sg13g2_decap_8
X_13296_ VGND VPWR net1678 _07008_ _00838_ _07009_ sg13g2_a21oi_1
X_12316_ _06162_ _06080_ _06161_ VPWR VGND sg13g2_nand2_1
XFILLER_54_7 VPWR VGND sg13g2_decap_8
XFILLER_5_374 VPWR VGND sg13g2_fill_1
XFILLER_114_228 VPWR VGND sg13g2_decap_8
X_12247_ _06093_ _06089_ _06092_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_21 VPWR VGND sg13g2_decap_8
XFILLER_111_957 VPWR VGND sg13g2_decap_8
XFILLER_96_624 VPWR VGND sg13g2_fill_1
X_12178_ VPWR _06024_ _06023_ VGND sg13g2_inv_1
XFILLER_1_580 VPWR VGND sg13g2_decap_8
X_11129_ _05099_ net1698 _05085_ VPWR VGND sg13g2_nand2_1
XFILLER_3_98 VPWR VGND sg13g2_decap_8
XFILLER_110_489 VPWR VGND sg13g2_decap_8
XFILLER_110_478 VPWR VGND sg13g2_fill_1
XFILLER_97_1012 VPWR VGND sg13g2_fill_2
XFILLER_76_370 VPWR VGND sg13g2_fill_1
X_14819_ _00620_ VGND VPWR _01343_ acc_sum.add_renorm0.mantisa\[8\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_1
XFILLER_91_340 VPWR VGND sg13g2_decap_8
XFILLER_24_418 VPWR VGND sg13g2_decap_8
XFILLER_45_790 VPWR VGND sg13g2_decap_8
X_08340_ sipo.word\[2\] sipo.word\[1\] sipo.word\[3\] _02585_ VPWR VGND sipo.word\[0\]
+ sg13g2_nand4_1
XFILLER_33_974 VPWR VGND sg13g2_decap_8
XFILLER_60_782 VPWR VGND sg13g2_decap_8
X_08271_ _02519_ VPWR _02520_ VGND _02467_ _02345_ sg13g2_o21ai_1
XFILLER_32_473 VPWR VGND sg13g2_decap_8
X_07222_ _01594_ acc_sub.op_sign_logic0.s_b acc_sub.op_sign_logic0.add_sub VPWR VGND
+ sg13g2_xnor2_1
XFILLER_80_0 VPWR VGND sg13g2_decap_4
X_07153_ VPWR _01525_ acc_sub.op_sign_logic0.mantisa_b\[6\] VGND sg13g2_inv_1
XFILLER_118_556 VPWR VGND sg13g2_fill_2
XFILLER_9_691 VPWR VGND sg13g2_fill_1
XFILLER_105_206 VPWR VGND sg13g2_fill_2
XFILLER_114_762 VPWR VGND sg13g2_decap_8
Xclkbuf_5_28__f_clk clknet_4_14_0_clk clknet_5_28__leaf_clk VPWR VGND sg13g2_buf_8
Xfanout103 net104 net103 VPWR VGND sg13g2_buf_2
XFILLER_99_462 VPWR VGND sg13g2_decap_8
XFILLER_99_451 VPWR VGND sg13g2_decap_8
Xfanout136 net140 net136 VPWR VGND sg13g2_buf_2
XFILLER_101_423 VPWR VGND sg13g2_decap_8
XFILLER_87_635 VPWR VGND sg13g2_decap_8
Xfanout125 net127 net125 VPWR VGND sg13g2_buf_2
Xfanout114 net116 net114 VPWR VGND sg13g2_buf_2
XFILLER_102_979 VPWR VGND sg13g2_decap_8
XFILLER_75_819 VPWR VGND sg13g2_decap_8
XFILLER_75_808 VPWR VGND sg13g2_fill_1
XFILLER_41_1000 VPWR VGND sg13g2_decap_8
X_07986_ _02256_ fp16_sum_pipe.exp_mant_logic0.a\[9\] _02250_ fp16_sum_pipe.seg_reg0.q\[24\]
+ net1775 VPWR VGND sg13g2_a22oi_1
XFILLER_74_318 VPWR VGND sg13g2_decap_8
XFILLER_110_990 VPWR VGND sg13g2_decap_8
X_09656_ _03772_ VPWR _03773_ VGND _03732_ _03726_ sg13g2_o21ai_1
XFILLER_83_852 VPWR VGND sg13g2_decap_8
XFILLER_28_768 VPWR VGND sg13g2_decap_4
XFILLER_103_66 VPWR VGND sg13g2_fill_1
X_08607_ acc_sum.op_sign_logic0.mantisa_a\[5\] acc_sum.op_sign_logic0.mantisa_b\[5\]
+ net1739 _02830_ VPWR VGND sg13g2_nand3_1
XFILLER_83_874 VPWR VGND sg13g2_fill_2
XFILLER_55_576 VPWR VGND sg13g2_decap_8
X_09587_ VPWR _03704_ _03703_ VGND sg13g2_inv_1
XFILLER_55_598 VPWR VGND sg13g2_fill_1
XFILLER_42_226 VPWR VGND sg13g2_decap_4
X_08538_ _02762_ _02761_ acc_sum.op_sign_logic0.mantisa_a\[0\] VPWR VGND sg13g2_nand2_1
XFILLER_42_248 VPWR VGND sg13g2_fill_2
XFILLER_24_974 VPWR VGND sg13g2_decap_8
X_08469_ _02701_ fpdiv.divider0.remainder_reg\[10\] net1708 _01756_ fpdiv.divider0.dividend\[10\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_10_112 VPWR VGND sg13g2_decap_8
X_10500_ VGND VPWR _04543_ net1848 _01168_ _04544_ sg13g2_a21oi_1
XFILLER_11_646 VPWR VGND sg13g2_decap_8
XFILLER_11_657 VPWR VGND sg13g2_fill_1
X_11480_ _05392_ VPWR _01036_ VGND fpdiv.reg1en.d\[0\] _05391_ sg13g2_o21ai_1
XFILLER_7_628 VPWR VGND sg13g2_fill_1
XFILLER_6_105 VPWR VGND sg13g2_decap_8
X_10431_ VPWR _04480_ _04479_ VGND sg13g2_inv_1
XFILLER_12_63 VPWR VGND sg13g2_decap_8
X_13150_ _00871_ _06896_ _06889_ VPWR VGND sg13g2_nand2_1
X_10362_ _04412_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[1\] VPWR VGND fp16_sum_pipe.op_sign_logic0.mantisa_b\[1\]
+ sg13g2_nand2b_2
XFILLER_124_548 VPWR VGND sg13g2_decap_4
X_13081_ _06846_ _06845_ _06813_ VPWR VGND sg13g2_nand2_1
X_12101_ _05947_ _05945_ _05946_ VPWR VGND sg13g2_nand2_1
X_10293_ _04298_ _04189_ _04361_ VPWR VGND sg13g2_nor2_1
X_12032_ _05876_ _05840_ _05879_ VPWR VGND sg13g2_nor2_1
XFILLER_3_889 VPWR VGND sg13g2_decap_8
XFILLER_2_388 VPWR VGND sg13g2_decap_8
XFILLER_120_743 VPWR VGND sg13g2_decap_8
XFILLER_104_294 VPWR VGND sg13g2_decap_8
XFILLER_78_679 VPWR VGND sg13g2_fill_2
XFILLER_78_668 VPWR VGND sg13g2_fill_1
X_13983_ VPWR _00534_ net13 VGND sg13g2_inv_1
XFILLER_101_990 VPWR VGND sg13g2_decap_8
XFILLER_93_649 VPWR VGND sg13g2_decap_8
XFILLER_74_841 VPWR VGND sg13g2_decap_8
XFILLER_58_392 VPWR VGND sg13g2_fill_1
X_12934_ _06707_ net1910 fp16_res_pipe.y\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_61_502 VPWR VGND sg13g2_decap_8
XFILLER_46_565 VPWR VGND sg13g2_decap_4
XFILLER_73_373 VPWR VGND sg13g2_fill_2
X_12865_ VPWR _06644_ fpmul.reg_p_out\[9\] VGND sg13g2_inv_1
X_12796_ _00020_ net1730 net1701 _06580_ VPWR VGND sg13g2_nand3_1
X_14604_ _00405_ VGND VPWR _01136_ fp16_res_pipe.y\[15\] clknet_leaf_128_clk sg13g2_dfrbpq_2
X_11816_ _05717_ _05573_ add_result\[11\] VPWR VGND sg13g2_nand2_1
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_18_1013 VPWR VGND sg13g2_fill_1
X_14535_ _00336_ VGND VPWR _01071_ fpdiv.div_out\[10\] clknet_leaf_76_clk sg13g2_dfrbpq_1
XFILLER_42_760 VPWR VGND sg13g2_decap_4
X_11747_ net1839 fp16_sum_pipe.add_renorm0.exp\[7\] _05651_ VPWR VGND sg13g2_nor2_1
XFILLER_14_451 VPWR VGND sg13g2_decap_8
XFILLER_30_955 VPWR VGND sg13g2_decap_8
X_14466_ _00267_ VGND VPWR _01005_ fpmul.seg_reg0.q\[51\] clknet_leaf_93_clk sg13g2_dfrbpq_1
X_11678_ VPWR _05582_ _05581_ VGND sg13g2_inv_1
X_14397_ _00198_ VGND VPWR _00936_ div_result\[10\] clknet_leaf_90_clk sg13g2_dfrbpq_1
X_13417_ _07087_ VPWR _00795_ VGND _07042_ net1722 sg13g2_o21ai_1
X_10629_ _04641_ VPWR _04642_ VGND fp16_res_pipe.add_renorm0.mantisa\[3\] _04640_
+ sg13g2_o21ai_1
XFILLER_127_364 VPWR VGND sg13g2_decap_8
Xplace1806 net1805 net1806 VPWR VGND sg13g2_buf_1
Xplace1817 net1816 net1817 VPWR VGND sg13g2_buf_2
X_13348_ _07048_ net1723 fp16_res_pipe.x2\[6\] VPWR VGND sg13g2_nand2_1
Xplace1828 fp16_res_pipe.exp_mant_logic0.a\[5\] net1828 VPWR VGND sg13g2_buf_2
Xplace1839 net1838 net1839 VPWR VGND sg13g2_buf_2
X_13279_ _03966_ _02573_ _06996_ VPWR VGND sg13g2_nor2_1
XFILLER_69_602 VPWR VGND sg13g2_decap_4
XFILLER_64_1000 VPWR VGND sg13g2_decap_8
XFILLER_123_581 VPWR VGND sg13g2_decap_8
XFILLER_96_421 VPWR VGND sg13g2_fill_1
XFILLER_69_635 VPWR VGND sg13g2_decap_8
XFILLER_69_613 VPWR VGND sg13g2_fill_2
XFILLER_111_754 VPWR VGND sg13g2_decap_8
XFILLER_110_242 VPWR VGND sg13g2_decap_8
X_07840_ _02136_ _02129_ _02135_ VPWR VGND sg13g2_nand2_1
XFILLER_97_977 VPWR VGND sg13g2_decap_8
XFILLER_96_432 VPWR VGND sg13g2_decap_8
X_07771_ _01418_ _02071_ _02072_ VPWR VGND sg13g2_nand2_1
XFILLER_96_465 VPWR VGND sg13g2_fill_2
XFILLER_84_616 VPWR VGND sg13g2_fill_2
XFILLER_56_329 VPWR VGND sg13g2_decap_8
X_09510_ _03619_ _03625_ _03627_ VPWR VGND sg13g2_nor2_1
XFILLER_49_370 VPWR VGND sg13g2_decap_8
XFILLER_37_510 VPWR VGND sg13g2_decap_8
XFILLER_25_705 VPWR VGND sg13g2_decap_8
XFILLER_65_896 VPWR VGND sg13g2_decap_4
X_09441_ _03579_ VPWR _01262_ VGND net1834 _03578_ sg13g2_o21ai_1
XFILLER_25_738 VPWR VGND sg13g2_decap_4
X_09372_ VGND VPWR _03430_ _03388_ _03521_ _03385_ sg13g2_a21oi_1
X_08323_ _02568_ _02567_ state\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_33_782 VPWR VGND sg13g2_decap_8
XFILLER_60_590 VPWR VGND sg13g2_fill_2
XFILLER_21_966 VPWR VGND sg13g2_decap_8
XFILLER_32_281 VPWR VGND sg13g2_fill_1
XFILLER_119_821 VPWR VGND sg13g2_decap_8
X_08254_ _02505_ fp16_sum_pipe.exp_mant_logic0.b\[2\] _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[5\]
+ net1777 VPWR VGND sg13g2_a22oi_1
XFILLER_20_454 VPWR VGND sg13g2_decap_4
X_07205_ _01576_ VPWR _01577_ VGND _01530_ _01575_ sg13g2_o21ai_1
X_08185_ _02443_ _02442_ net1639 VPWR VGND sg13g2_nand2_1
XFILLER_119_898 VPWR VGND sg13g2_decap_8
X_07136_ VPWR _01508_ _01507_ VGND sg13g2_inv_1
XFILLER_118_397 VPWR VGND sg13g2_decap_8
XFILLER_106_526 VPWR VGND sg13g2_decap_8
XFILLER_3_119 VPWR VGND sg13g2_decap_8
XFILLER_88_900 VPWR VGND sg13g2_fill_1
XFILLER_59_112 VPWR VGND sg13g2_decap_8
XFILLER_58_37 VPWR VGND sg13g2_fill_2
XFILLER_58_26 VPWR VGND sg13g2_fill_2
XFILLER_58_59 VPWR VGND sg13g2_fill_1
XFILLER_114_21 VPWR VGND sg13g2_decap_8
XFILLER_88_988 VPWR VGND sg13g2_decap_8
XFILLER_68_690 VPWR VGND sg13g2_decap_8
X_07969_ _02242_ VPWR _02243_ VGND fp16_sum_pipe.exp_mant_logic0.b\[13\] _02241_ sg13g2_o21ai_1
XFILLER_114_98 VPWR VGND sg13g2_decap_8
XFILLER_74_159 VPWR VGND sg13g2_decap_8
XFILLER_56_863 VPWR VGND sg13g2_decap_8
X_10980_ _04976_ fp16_res_pipe.x2\[14\] net1926 VPWR VGND sg13g2_nand2_1
X_09639_ net1804 VPWR _03756_ VGND _03751_ _03755_ sg13g2_o21ai_1
XFILLER_70_321 VPWR VGND sg13g2_decap_8
XFILLER_16_749 VPWR VGND sg13g2_fill_2
X_12650_ VPWR _06466_ _06465_ VGND sg13g2_inv_1
XFILLER_70_332 VPWR VGND sg13g2_fill_2
XFILLER_43_546 VPWR VGND sg13g2_decap_8
XFILLER_12_911 VPWR VGND sg13g2_decap_8
X_11601_ _05430_ _05462_ _05506_ VPWR VGND sg13g2_nor2_1
X_12581_ _06378_ _06381_ _06397_ VPWR VGND sg13g2_xor2_1
XFILLER_51_590 VPWR VGND sg13g2_fill_1
X_14320_ _00121_ VGND VPWR _00863_ sipo.word\[8\] clknet_leaf_12_clk sg13g2_dfrbpq_2
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_12_988 VPWR VGND sg13g2_decap_8
X_11532_ fp16_sum_pipe.add_renorm0.mantisa\[4\] fp16_sum_pipe.add_renorm0.mantisa\[3\]
+ fp16_sum_pipe.add_renorm0.mantisa\[5\] _05437_ VPWR VGND sg13g2_nand3_1
X_11463_ _05384_ VPWR _01045_ VGND net1947 _02722_ sg13g2_o21ai_1
XFILLER_87_1000 VPWR VGND sg13g2_decap_8
X_14251_ _00052_ VGND VPWR _00802_ acc_sub.x2\[0\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_7_447 VPWR VGND sg13g2_decap_4
XFILLER_23_84 VPWR VGND sg13g2_decap_8
XFILLER_125_802 VPWR VGND sg13g2_decap_8
XFILLER_124_301 VPWR VGND sg13g2_decap_8
X_14182_ VPWR _00733_ net116 VGND sg13g2_inv_1
X_13202_ _06936_ net1714 sipo.word\[3\] VPWR VGND sg13g2_nand2_1
X_10414_ _04463_ VPWR _04464_ VGND fp16_sum_pipe.op_sign_logic0.s_a _04460_ sg13g2_o21ai_1
X_11394_ _05341_ net1718 fpdiv.div_out\[8\] VPWR VGND sg13g2_nand2_1
X_13133_ _06885_ _06573_ _06882_ VPWR VGND sg13g2_nand2_1
XFILLER_125_879 VPWR VGND sg13g2_decap_8
XFILLER_124_356 VPWR VGND sg13g2_fill_1
XFILLER_112_507 VPWR VGND sg13g2_decap_4
XFILLER_3_653 VPWR VGND sg13g2_decap_8
X_10345_ _04395_ _04393_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[9\] VPWR VGND sg13g2_nand2_1
X_13064_ _05815_ _05817_ _05809_ _06832_ VPWR VGND _05821_ sg13g2_nand4_1
X_10276_ _04346_ _04340_ _04345_ VPWR VGND sg13g2_nand2_1
XFILLER_94_903 VPWR VGND sg13g2_decap_4
X_12015_ _05866_ _05848_ _05847_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_196 VPWR VGND sg13g2_decap_8
Xclkbuf_5_11__f_clk clknet_4_5_0_clk clknet_5_11__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_78_476 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_39_819 VPWR VGND sg13g2_decap_8
XFILLER_94_947 VPWR VGND sg13g2_decap_8
XFILLER_93_435 VPWR VGND sg13g2_decap_8
XFILLER_66_649 VPWR VGND sg13g2_decap_8
XFILLER_59_690 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_65_159 VPWR VGND sg13g2_fill_2
XFILLER_46_340 VPWR VGND sg13g2_decap_8
XFILLER_19_543 VPWR VGND sg13g2_decap_8
X_13966_ VPWR _00517_ net7 VGND sg13g2_inv_1
X_12917_ _06692_ net1717 _00010_ VPWR VGND sg13g2_nand2_1
XFILLER_74_682 VPWR VGND sg13g2_decap_8
XFILLER_34_502 VPWR VGND sg13g2_fill_2
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_19_598 VPWR VGND sg13g2_fill_1
X_13897_ VPWR _00448_ net11 VGND sg13g2_inv_1
X_12848_ VGND VPWR net1935 add_result\[10\] _06628_ net1943 sg13g2_a21oi_1
XFILLER_62_899 VPWR VGND sg13g2_fill_2
XFILLER_61_387 VPWR VGND sg13g2_decap_8
XFILLER_22_719 VPWR VGND sg13g2_fill_1
X_12779_ VPWR _06564_ piso.tx_active VGND sg13g2_inv_1
XFILLER_9_42 VPWR VGND sg13g2_decap_8
XFILLER_14_292 VPWR VGND sg13g2_fill_1
X_14518_ _00319_ VGND VPWR _01054_ fpdiv.reg_a_out\[9\] clknet_leaf_54_clk sg13g2_dfrbpq_2
XFILLER_80_90 VPWR VGND sg13g2_decap_8
X_14449_ _00250_ VGND VPWR _00988_ fpmul.seg_reg0.q\[34\] clknet_leaf_97_clk sg13g2_dfrbpq_1
XFILLER_30_785 VPWR VGND sg13g2_fill_2
XFILLER_127_161 VPWR VGND sg13g2_decap_8
XFILLER_116_835 VPWR VGND sg13g2_decap_8
XFILLER_115_334 VPWR VGND sg13g2_decap_8
Xplace1636 _04272_ net1636 VPWR VGND sg13g2_buf_2
XFILLER_115_367 VPWR VGND sg13g2_fill_2
Xplace1669 _01844_ net1669 VPWR VGND sg13g2_buf_2
XFILLER_103_507 VPWR VGND sg13g2_decap_8
Xplace1647 _02692_ net1647 VPWR VGND sg13g2_buf_2
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_09990_ _04042_ VPWR _04078_ VGND _03996_ _04077_ sg13g2_o21ai_1
Xplace1658 _02347_ net1658 VPWR VGND sg13g2_buf_2
X_08941_ _03128_ _03010_ _02967_ VPWR VGND sg13g2_nand2_1
XFILLER_9_1011 VPWR VGND sg13g2_fill_2
X_08872_ VPWR _03059_ _03058_ VGND sg13g2_inv_1
X_07823_ _02120_ acc_sub.exp_mant_logic0.b\[1\] net1651 net1685 acc_sub.exp_mant_logic0.b\[0\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_85_936 VPWR VGND sg13g2_decap_8
XFILLER_38_841 VPWR VGND sg13g2_decap_8
X_07754_ _02055_ _02056_ _02054_ _02058_ VPWR VGND _02057_ sg13g2_nand4_1
XFILLER_84_468 VPWR VGND sg13g2_fill_2
XFILLER_84_457 VPWR VGND sg13g2_decap_8
X_07685_ _01994_ acc_sub.exp_mant_logic0.a\[2\] _01923_ _01871_ acc_sub.exp_mant_logic0.a\[1\]
+ VPWR VGND sg13g2_a22oi_1
Xclkbuf_leaf_91_clk clknet_5_13__leaf_clk clknet_leaf_91_clk VPWR VGND sg13g2_buf_8
XFILLER_53_866 VPWR VGND sg13g2_decap_8
XFILLER_53_844 VPWR VGND sg13g2_fill_1
XFILLER_44_28 VPWR VGND sg13g2_decap_8
X_09424_ _03567_ net1675 _03449_ VPWR VGND sg13g2_nand2_1
X_09355_ VGND VPWR _03433_ _03436_ _03506_ _03371_ sg13g2_a21oi_1
X_08306_ _02552_ net1657 fp16_sum_pipe.exp_mant_logic0.b\[2\] VPWR VGND sg13g2_nand2_1
X_09286_ _03369_ _03439_ _03440_ VPWR VGND sg13g2_nor2_1
XFILLER_121_7 VPWR VGND sg13g2_decap_8
X_08237_ _02490_ fp16_sum_pipe.exp_mant_logic0.b\[4\] _02246_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[7\]
+ net1778 VPWR VGND sg13g2_a22oi_1
XFILLER_109_21 VPWR VGND sg13g2_decap_8
XFILLER_4_406 VPWR VGND sg13g2_decap_8
XFILLER_118_161 VPWR VGND sg13g2_decap_8
XFILLER_69_14 VPWR VGND sg13g2_decap_8
X_08168_ _02427_ _02307_ _02426_ VPWR VGND sg13g2_nand2_2
XFILLER_122_805 VPWR VGND sg13g2_decap_8
X_07119_ VPWR _01492_ acc_sub.reg2en.q\[0\] VGND sg13g2_inv_1
XFILLER_69_25 VPWR VGND sg13g2_decap_8
X_08099_ _02363_ fp16_sum_pipe.exp_mant_logic0.a\[6\] net1659 net1691 fp16_sum_pipe.exp_mant_logic0.a\[4\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_106_389 VPWR VGND sg13g2_decap_8
XFILLER_79_207 VPWR VGND sg13g2_decap_4
XFILLER_69_69 VPWR VGND sg13g2_decap_8
X_10130_ _04211_ VPWR _04212_ VGND _03615_ _04124_ sg13g2_o21ai_1
XFILLER_125_42 VPWR VGND sg13g2_decap_8
XFILLER_88_730 VPWR VGND sg13g2_decap_4
X_10061_ _04133_ _04136_ _04148_ _04149_ VPWR VGND sg13g2_nor3_1
XFILLER_88_796 VPWR VGND sg13g2_decap_8
XFILLER_85_24 VPWR VGND sg13g2_decap_4
XFILLER_87_284 VPWR VGND sg13g2_decap_8
XFILLER_76_969 VPWR VGND sg13g2_decap_8
XFILLER_85_79 VPWR VGND sg13g2_fill_1
X_13820_ VPWR _00371_ net52 VGND sg13g2_inv_1
XFILLER_28_351 VPWR VGND sg13g2_fill_1
XFILLER_84_980 VPWR VGND sg13g2_decap_8
X_13751_ VPWR _00302_ net114 VGND sg13g2_inv_1
XFILLER_62_118 VPWR VGND sg13g2_fill_2
XFILLER_55_170 VPWR VGND sg13g2_decap_8
X_10963_ _04967_ VPWR _01128_ VGND _04966_ _04771_ sg13g2_o21ai_1
XFILLER_28_362 VPWR VGND sg13g2_decap_8
X_12702_ _06510_ div_result\[6\] VPWR VGND sg13g2_inv_2
Xclkbuf_leaf_82_clk clknet_5_24__leaf_clk clknet_leaf_82_clk VPWR VGND sg13g2_buf_8
XFILLER_55_181 VPWR VGND sg13g2_fill_1
XFILLER_16_535 VPWR VGND sg13g2_decap_4
XFILLER_70_151 VPWR VGND sg13g2_decap_4
X_13682_ VPWR _00233_ net69 VGND sg13g2_inv_1
X_10894_ _04903_ _04791_ _04904_ VPWR VGND sg13g2_nor2b_1
X_12633_ _06440_ _06448_ _06449_ VPWR VGND sg13g2_nor2_1
X_12564_ _06380_ fpdiv.reg_a_out\[9\] fpdiv.reg_b_out\[9\] VPWR VGND sg13g2_xnor2_1
XFILLER_8_712 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_decap_8
X_14303_ _00104_ VGND VPWR _00847_ acc\[13\] clknet_leaf_23_clk sg13g2_dfrbpq_2
XFILLER_11_273 VPWR VGND sg13g2_decap_8
XFILLER_11_284 VPWR VGND sg13g2_fill_1
X_11515_ _05420_ net1841 fp16_sum_pipe.add_renorm0.mantisa\[7\] VPWR VGND sg13g2_nand2_1
X_12495_ _06233_ _06238_ _06330_ VPWR VGND sg13g2_nor2_1
X_14234_ _00035_ VGND VPWR _00785_ sipo.shift_reg\[15\] clknet_leaf_7_clk sg13g2_dfrbpq_1
XFILLER_7_233 VPWR VGND sg13g2_decap_8
X_11446_ _05373_ VPWR _01051_ VGND net1947 _05372_ sg13g2_o21ai_1
XFILLER_7_277 VPWR VGND sg13g2_fill_1
XFILLER_113_816 VPWR VGND sg13g2_decap_8
X_14165_ VPWR _00716_ net103 VGND sg13g2_inv_1
X_11377_ _05324_ _05327_ _05328_ VPWR VGND _05320_ sg13g2_nand3b_1
XFILLER_4_951 VPWR VGND sg13g2_decap_8
XFILLER_124_175 VPWR VGND sg13g2_decap_8
XFILLER_112_315 VPWR VGND sg13g2_decap_8
X_13116_ _06872_ VPWR _00881_ VGND net1862 _06710_ sg13g2_o21ai_1
X_14096_ VPWR _00647_ net41 VGND sg13g2_inv_1
X_10328_ _04381_ VPWR _01177_ VGND net1921 _04298_ sg13g2_o21ai_1
XFILLER_98_549 VPWR VGND sg13g2_decap_8
X_13047_ VPWR _06815_ _06814_ VGND sg13g2_inv_1
XFILLER_3_483 VPWR VGND sg13g2_decap_8
XFILLER_121_882 VPWR VGND sg13g2_decap_8
XFILLER_66_402 VPWR VGND sg13g2_decap_8
X_10259_ _04330_ net1644 fp16_res_pipe.exp_mant_logic0.b\[1\] VPWR VGND sg13g2_nand2_1
XFILLER_38_126 VPWR VGND sg13g2_decap_8
XFILLER_94_766 VPWR VGND sg13g2_decap_8
XFILLER_93_243 VPWR VGND sg13g2_decap_8
XFILLER_66_479 VPWR VGND sg13g2_decap_8
XFILLER_93_276 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_73_clk clknet_5_31__leaf_clk clknet_leaf_73_clk VPWR VGND sg13g2_buf_8
X_13949_ VPWR _00500_ net97 VGND sg13g2_inv_1
X_07470_ _01787_ _01792_ _01793_ VPWR VGND sg13g2_nor2_1
XFILLER_62_674 VPWR VGND sg13g2_decap_8
XFILLER_61_140 VPWR VGND sg13g2_decap_8
XFILLER_22_516 VPWR VGND sg13g2_fill_1
XFILLER_34_387 VPWR VGND sg13g2_fill_1
X_09140_ VGND VPWR _03316_ _03318_ _03319_ _03136_ sg13g2_a21oi_1
X_09071_ _03237_ _03239_ _03256_ VPWR VGND sg13g2_xor2_1
X_08022_ VGND VPWR _02233_ _02196_ _02288_ _02193_ sg13g2_a21oi_1
XFILLER_116_632 VPWR VGND sg13g2_decap_4
Xfanout5 net6 net5 VPWR VGND sg13g2_buf_2
XFILLER_115_175 VPWR VGND sg13g2_decap_8
X_09973_ _04063_ _04064_ _04062_ _01215_ VPWR VGND sg13g2_nand3_1
X_08924_ _03110_ _03067_ _03111_ VPWR VGND sg13g2_xor2_1
XFILLER_39_28 VPWR VGND sg13g2_decap_8
XFILLER_69_262 VPWR VGND sg13g2_decap_4
XFILLER_69_240 VPWR VGND sg13g2_fill_1
XFILLER_58_925 VPWR VGND sg13g2_decap_8
XFILLER_58_903 VPWR VGND sg13g2_decap_8
XFILLER_57_402 VPWR VGND sg13g2_decap_8
X_08855_ _03042_ _03036_ _03038_ _03041_ VPWR VGND sg13g2_and3_2
XFILLER_85_733 VPWR VGND sg13g2_decap_8
X_08786_ VPWR _02973_ _02971_ VGND sg13g2_inv_1
X_07806_ _02104_ _02102_ _02103_ VPWR VGND sg13g2_nand2_1
XFILLER_85_755 VPWR VGND sg13g2_fill_2
XFILLER_84_254 VPWR VGND sg13g2_decap_8
XFILLER_29_148 VPWR VGND sg13g2_decap_8
X_07737_ VPWR _02042_ acc_sub.op_sign_logic0.mantisa_a\[0\] VGND sg13g2_inv_1
XFILLER_72_416 VPWR VGND sg13g2_decap_8
XFILLER_55_49 VPWR VGND sg13g2_decap_8
XFILLER_38_671 VPWR VGND sg13g2_decap_8
XFILLER_81_950 VPWR VGND sg13g2_decap_8
X_07668_ _01868_ _01977_ _01978_ VPWR VGND sg13g2_nor2_1
XFILLER_80_471 VPWR VGND sg13g2_decap_8
XFILLER_53_685 VPWR VGND sg13g2_fill_2
XFILLER_13_516 VPWR VGND sg13g2_decap_4
XFILLER_111_77 VPWR VGND sg13g2_decap_8
X_07599_ _01912_ _01810_ _01913_ VPWR VGND sg13g2_xor2_1
X_09407_ _03551_ VPWR _03552_ VGND net1675 _03550_ sg13g2_o21ai_1
XFILLER_40_368 VPWR VGND sg13g2_decap_8
X_09338_ VGND VPWR _03489_ _03407_ _03490_ _03404_ sg13g2_a21oi_1
X_11300_ _05259_ net1811 net1681 acc_sum.op_sign_logic0.mantisa_b\[9\] net1762 VPWR
+ VGND sg13g2_a22oi_1
X_09269_ VPWR _03423_ fp16_res_pipe.op_sign_logic0.mantisa_a\[4\] VGND sg13g2_inv_1
XFILLER_126_429 VPWR VGND sg13g2_fill_1
X_12280_ _06126_ _06125_ _06116_ VPWR VGND sg13g2_nand2_1
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_106_142 VPWR VGND sg13g2_fill_1
XFILLER_106_131 VPWR VGND sg13g2_fill_2
X_11231_ _02953_ _05148_ _05196_ VPWR VGND sg13g2_nor2_1
XFILLER_5_759 VPWR VGND sg13g2_decap_8
X_11162_ _05119_ _05116_ _05131_ VPWR VGND sg13g2_nor2_1
XFILLER_20_63 VPWR VGND sg13g2_decap_8
XFILLER_121_112 VPWR VGND sg13g2_decap_8
X_10113_ net1746 _04128_ _04195_ _04196_ VPWR VGND sg13g2_nand3_1
XFILLER_110_808 VPWR VGND sg13g2_decap_8
XFILLER_96_56 VPWR VGND sg13g2_decap_8
X_11093_ _05066_ net1760 acc_sum.seg_reg0.q\[23\] VPWR VGND sg13g2_nand2_1
XFILLER_0_442 VPWR VGND sg13g2_decap_8
XFILLER_1_976 VPWR VGND sg13g2_decap_8
XFILLER_121_189 VPWR VGND sg13g2_decap_8
X_14921_ _00722_ VGND VPWR _01441_ acc_sub.op_sign_logic0.s_b clknet_leaf_43_clk sg13g2_dfrbpq_2
XFILLER_88_593 VPWR VGND sg13g2_fill_1
XFILLER_76_733 VPWR VGND sg13g2_decap_8
XFILLER_76_722 VPWR VGND sg13g2_decap_4
XFILLER_49_958 VPWR VGND sg13g2_decap_8
XFILLER_48_435 VPWR VGND sg13g2_decap_4
XFILLER_64_906 VPWR VGND sg13g2_fill_2
X_14852_ _00653_ VGND VPWR _01376_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[3\] clknet_leaf_112_clk
+ sg13g2_dfrbpq_1
XFILLER_29_72 VPWR VGND sg13g2_fill_1
X_13803_ VPWR _00354_ net81 VGND sg13g2_inv_1
XFILLER_17_800 VPWR VGND sg13g2_fill_2
X_14783_ _00584_ VGND VPWR _01307_ acc_sub.y\[12\] clknet_leaf_39_clk sg13g2_dfrbpq_1
XFILLER_90_246 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_55_clk clknet_5_19__leaf_clk clknet_leaf_55_clk VPWR VGND sg13g2_buf_8
XFILLER_56_490 VPWR VGND sg13g2_decap_8
X_11995_ _05849_ _05847_ _05848_ VPWR VGND sg13g2_nand2_1
XFILLER_16_310 VPWR VGND sg13g2_decap_8
XFILLER_29_693 VPWR VGND sg13g2_fill_2
XFILLER_90_268 VPWR VGND sg13g2_fill_1
XFILLER_90_257 VPWR VGND sg13g2_decap_8
X_13734_ VPWR _00285_ net63 VGND sg13g2_inv_1
XFILLER_43_140 VPWR VGND sg13g2_decap_8
XFILLER_17_877 VPWR VGND sg13g2_decap_8
X_10946_ _04737_ _04951_ _04952_ VPWR VGND _04844_ sg13g2_nand3b_1
XFILLER_32_825 VPWR VGND sg13g2_fill_1
X_13665_ VPWR _00216_ net36 VGND sg13g2_inv_1
XFILLER_43_162 VPWR VGND sg13g2_decap_8
X_10877_ VPWR _04888_ _04887_ VGND sg13g2_inv_1
XFILLER_31_313 VPWR VGND sg13g2_decap_8
X_12616_ _06427_ _06431_ _06432_ VPWR VGND sg13g2_nor2_1
XFILLER_31_346 VPWR VGND sg13g2_fill_2
XFILLER_118_908 VPWR VGND sg13g2_decap_8
XFILLER_84_7 VPWR VGND sg13g2_fill_2
X_13596_ VPWR _00147_ net110 VGND sg13g2_inv_1
XFILLER_40_880 VPWR VGND sg13g2_decap_8
X_12547_ fpdiv.reg_b_out\[13\] fpdiv.reg_b_out\[12\] fpdiv.reg_b_out\[11\] fpdiv.reg_b_out\[10\]
+ _06364_ VPWR VGND sg13g2_nor4_1
XFILLER_61_81 VPWR VGND sg13g2_decap_8
X_12478_ net1872 fpmul.seg_reg0.q\[9\] _06318_ VPWR VGND sg13g2_nor2_1
XFILLER_6_21 VPWR VGND sg13g2_decap_8
XFILLER_126_974 VPWR VGND sg13g2_decap_8
X_14217_ VPWR _00768_ net133 VGND sg13g2_inv_1
X_11429_ _05362_ VPWR _01057_ VGND net1938 _05361_ sg13g2_o21ai_1
X_14148_ VPWR _00699_ net134 VGND sg13g2_inv_1
XFILLER_6_98 VPWR VGND sg13g2_decap_8
Xclkbuf_5_9__f_clk clknet_4_4_0_clk clknet_5_9__leaf_clk VPWR VGND sg13g2_buf_8
X_14079_ VPWR _00630_ net137 VGND sg13g2_inv_1
XFILLER_100_307 VPWR VGND sg13g2_decap_8
XFILLER_79_560 VPWR VGND sg13g2_decap_8
XFILLER_67_700 VPWR VGND sg13g2_decap_8
XFILLER_112_178 VPWR VGND sg13g2_fill_1
X_08640_ VGND VPWR _02860_ net1818 _01345_ _02861_ sg13g2_a21oi_1
XFILLER_94_585 VPWR VGND sg13g2_decap_4
XFILLER_27_619 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_46_clk clknet_5_22__leaf_clk clknet_leaf_46_clk VPWR VGND sg13g2_buf_8
X_08571_ VPWR _02795_ acc_sum.op_sign_logic0.mantisa_a\[10\] VGND sg13g2_inv_1
XFILLER_19_170 VPWR VGND sg13g2_fill_1
XFILLER_26_129 VPWR VGND sg13g2_fill_2
X_07522_ VPWR _01843_ net1686 VGND sg13g2_inv_1
XFILLER_62_460 VPWR VGND sg13g2_decap_4
XFILLER_35_663 VPWR VGND sg13g2_decap_8
XFILLER_34_140 VPWR VGND sg13g2_decap_8
X_07453_ VGND VPWR net1796 _01776_ _01441_ _01777_ sg13g2_a21oi_1
XFILLER_62_493 VPWR VGND sg13g2_decap_8
XFILLER_34_184 VPWR VGND sg13g2_fill_2
XFILLER_22_302 VPWR VGND sg13g2_fill_2
XFILLER_22_324 VPWR VGND sg13g2_decap_4
XFILLER_23_836 VPWR VGND sg13g2_decap_8
XFILLER_22_335 VPWR VGND sg13g2_decap_8
X_09123_ _03301_ _03303_ _03135_ _03304_ VPWR VGND sg13g2_nand3_1
X_07384_ _01731_ acc_sub.exp_mant_logic0.a\[11\] VPWR VGND sg13g2_inv_2
XFILLER_31_880 VPWR VGND sg13g2_fill_2
X_09054_ _03237_ _03239_ _03240_ VPWR VGND sg13g2_nor2b_1
XFILLER_108_418 VPWR VGND sg13g2_decap_8
XFILLER_117_963 VPWR VGND sg13g2_decap_8
X_08005_ _02263_ _02265_ _02266_ _02272_ VGND VPWR _02271_ sg13g2_nor4_2
XFILLER_103_101 VPWR VGND sg13g2_decap_8
XFILLER_103_167 VPWR VGND sg13g2_decap_8
X_09956_ _04051_ net1689 VPWR VGND sg13g2_inv_2
X_08907_ _03016_ _03093_ _03094_ VPWR VGND sg13g2_nor2b_2
X_09887_ net1831 fp16_res_pipe.op_sign_logic0.s_b _03986_ VPWR VGND sg13g2_nor2_1
X_08838_ VPWR _03025_ acc_sub.add_renorm0.mantisa\[3\] VGND sg13g2_inv_1
XFILLER_122_21 VPWR VGND sg13g2_decap_8
XFILLER_85_574 VPWR VGND sg13g2_decap_8
XFILLER_73_736 VPWR VGND sg13g2_decap_8
XFILLER_46_939 VPWR VGND sg13g2_fill_1
XFILLER_39_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_37_clk clknet_5_21__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
X_08769_ _02959_ acc_sum.exp_mant_logic0.a\[2\] VPWR VGND sg13g2_inv_2
XFILLER_122_98 VPWR VGND sg13g2_decap_8
XFILLER_60_408 VPWR VGND sg13g2_fill_1
X_11780_ _05682_ _05648_ _05681_ _05683_ VPWR VGND sg13g2_nand3_1
XFILLER_25_151 VPWR VGND sg13g2_fill_1
X_10800_ VPWR _04812_ _04811_ VGND sg13g2_inv_1
XFILLER_82_69 VPWR VGND sg13g2_decap_8
XFILLER_14_825 VPWR VGND sg13g2_decap_8
X_10731_ _04741_ _04743_ _04744_ VPWR VGND sg13g2_nor2_1
XFILLER_26_685 VPWR VGND sg13g2_fill_1
X_13450_ _07104_ VPWR _00779_ VGND _06923_ net1754 sg13g2_o21ai_1
XFILLER_15_63 VPWR VGND sg13g2_decap_4
X_12401_ _06210_ _06246_ _06247_ VPWR VGND sg13g2_nor2_1
XFILLER_51_1013 VPWR VGND sg13g2_fill_1
XFILLER_41_688 VPWR VGND sg13g2_decap_4
XFILLER_40_154 VPWR VGND sg13g2_decap_8
X_10662_ _04675_ fp16_res_pipe.add_renorm0.mantisa\[6\] _04645_ VPWR VGND sg13g2_xnor2_1
X_13381_ _07067_ net1695 sipo.word\[8\] VPWR VGND sg13g2_nand2_1
X_10593_ _04609_ VPWR _01140_ VGND net1934 _02268_ sg13g2_o21ai_1
XFILLER_22_891 VPWR VGND sg13g2_decap_8
XFILLER_108_930 VPWR VGND sg13g2_decap_8
X_12332_ VPWR _06178_ _06172_ VGND sg13g2_inv_1
XFILLER_126_259 VPWR VGND sg13g2_decap_8
XFILLER_110_0 VPWR VGND sg13g2_decap_8
X_12263_ _06079_ _06083_ _06109_ VPWR VGND sg13g2_nor2_1
XFILLER_5_534 VPWR VGND sg13g2_decap_8
XFILLER_31_95 VPWR VGND sg13g2_decap_4
XFILLER_123_911 VPWR VGND sg13g2_decap_8
X_14002_ VPWR _00553_ net78 VGND sg13g2_inv_1
X_11214_ _05112_ _05144_ _05180_ VPWR VGND sg13g2_nor2_1
X_12194_ _06040_ _06037_ _06039_ VPWR VGND sg13g2_nand2_1
XFILLER_123_988 VPWR VGND sg13g2_decap_8
XFILLER_110_605 VPWR VGND sg13g2_fill_1
XFILLER_95_305 VPWR VGND sg13g2_decap_8
X_11145_ _05114_ VPWR _05115_ VGND _05032_ net1698 sg13g2_o21ai_1
XFILLER_49_700 VPWR VGND sg13g2_fill_1
XFILLER_1_751 VPWR VGND sg13g2_decap_8
XFILLER_122_498 VPWR VGND sg13g2_decap_8
XFILLER_49_711 VPWR VGND sg13g2_decap_8
X_14904_ _00705_ VGND VPWR _01424_ acc_sub.op_sign_logic0.mantisa_a\[3\] clknet_leaf_62_clk
+ sg13g2_dfrbpq_2
XFILLER_88_390 VPWR VGND sg13g2_decap_8
XFILLER_49_744 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
X_10027_ VPWR _04115_ _04114_ VGND sg13g2_inv_1
XFILLER_49_799 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
X_14835_ _00636_ VGND VPWR _01359_ state\[1\] clknet_leaf_52_clk sg13g2_dfrbpq_2
Xclkbuf_leaf_28_clk clknet_5_16__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
X_14766_ _00567_ VGND VPWR _01290_ acc_sum.exp_mant_logic0.b\[11\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_11978_ _05832_ fpmul.reg_a_out\[9\] fpmul.reg_b_out\[9\] VPWR VGND sg13g2_nand2_1
XFILLER_51_408 VPWR VGND sg13g2_decap_8
X_13717_ VPWR _00268_ net58 VGND sg13g2_inv_1
X_10929_ _04873_ _04871_ _04937_ VPWR VGND sg13g2_nor2_1
X_14697_ _00498_ VGND VPWR _01225_ acc_sum.y\[0\] clknet_leaf_38_clk sg13g2_dfrbpq_1
XFILLER_60_953 VPWR VGND sg13g2_decap_8
XFILLER_31_132 VPWR VGND sg13g2_decap_4
XFILLER_82_4 VPWR VGND sg13g2_fill_1
X_13648_ VPWR _00199_ net108 VGND sg13g2_inv_1
XFILLER_31_165 VPWR VGND sg13g2_decap_8
X_13579_ VPWR _00130_ net21 VGND sg13g2_inv_1
XFILLER_13_891 VPWR VGND sg13g2_decap_8
XFILLER_117_259 VPWR VGND sg13g2_decap_8
XFILLER_126_771 VPWR VGND sg13g2_decap_8
XFILLER_114_944 VPWR VGND sg13g2_decap_8
XFILLER_113_421 VPWR VGND sg13g2_decap_4
XFILLER_113_432 VPWR VGND sg13g2_decap_4
XFILLER_99_644 VPWR VGND sg13g2_fill_1
XFILLER_98_110 VPWR VGND sg13g2_decap_8
X_09810_ _03663_ VPWR _03923_ VGND _03922_ _03910_ sg13g2_o21ai_1
XFILLER_87_806 VPWR VGND sg13g2_decap_8
X_09741_ VGND VPWR _03856_ _03857_ _03810_ _03828_ sg13g2_a21oi_2
XFILLER_98_176 VPWR VGND sg13g2_fill_1
X_09672_ acc_sum.add_renorm0.exp\[1\] acc_sum.add_renorm0.exp\[0\] acc_sum.add_renorm0.exp\[2\]
+ _03788_ VPWR VGND sg13g2_nand3_1
XFILLER_27_405 VPWR VGND sg13g2_fill_2
XFILLER_27_416 VPWR VGND sg13g2_fill_1
XFILLER_28_917 VPWR VGND sg13g2_decap_8
X_08623_ _02760_ VPWR _02845_ VGND _02841_ _02765_ sg13g2_o21ai_1
Xclkbuf_leaf_19_clk clknet_5_18__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_54_235 VPWR VGND sg13g2_fill_1
XFILLER_54_224 VPWR VGND sg13g2_decap_8
XFILLER_39_298 VPWR VGND sg13g2_decap_8
X_08554_ _02778_ _02776_ acc_sum.op_sign_logic0.mantisa_b\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_70_706 VPWR VGND sg13g2_decap_4
XFILLER_54_257 VPWR VGND sg13g2_fill_2
XFILLER_36_983 VPWR VGND sg13g2_decap_8
X_07505_ _01826_ VPWR _01827_ VGND _01814_ _01812_ sg13g2_o21ai_1
XFILLER_74_1013 VPWR VGND sg13g2_fill_1
XFILLER_51_931 VPWR VGND sg13g2_decap_4
XFILLER_35_460 VPWR VGND sg13g2_decap_8
X_08485_ _02714_ fpdiv.divider0.remainder_reg\[7\] net1708 net1748 fpdiv.divider0.dividend\[7\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_62_290 VPWR VGND sg13g2_decap_8
XFILLER_52_28 VPWR VGND sg13g2_decap_8
X_07436_ VGND VPWR _01766_ net1750 _01448_ _01767_ sg13g2_a21oi_1
XFILLER_22_176 VPWR VGND sg13g2_decap_4
XFILLER_23_677 VPWR VGND sg13g2_decap_8
X_07367_ _01720_ VPWR _01470_ VGND net1798 _01719_ sg13g2_o21ai_1
X_09106_ _03206_ _03205_ _03288_ VPWR VGND sg13g2_nor2_1
X_07298_ _01664_ net1667 _01629_ VPWR VGND sg13g2_nand2_1
X_09037_ VPWR _03223_ _03222_ VGND sg13g2_inv_1
XFILLER_108_237 VPWR VGND sg13g2_decap_4
XFILLER_117_760 VPWR VGND sg13g2_decap_8
XFILLER_117_21 VPWR VGND sg13g2_decap_8
XFILLER_105_944 VPWR VGND sg13g2_decap_8
XFILLER_104_443 VPWR VGND sg13g2_decap_8
XFILLER_81_1006 VPWR VGND sg13g2_decap_8
XFILLER_78_828 VPWR VGND sg13g2_fill_2
XFILLER_120_925 VPWR VGND sg13g2_decap_8
XFILLER_117_98 VPWR VGND sg13g2_decap_8
Xclkbuf_4_13_0_clk clknet_0_clk clknet_4_13_0_clk VPWR VGND sg13g2_buf_8
X_09939_ _04035_ _04034_ fp16_res_pipe.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_92_308 VPWR VGND sg13g2_fill_2
X_12950_ _06722_ _06721_ net1961 VPWR VGND sg13g2_nand2_1
XFILLER_93_35 VPWR VGND sg13g2_decap_8
X_12881_ _06659_ _06574_ _00013_ VPWR VGND sg13g2_nand2_1
XFILLER_73_533 VPWR VGND sg13g2_decap_8
X_11901_ fpmul.seg_reg0.q\[49\] fpmul.reg_a_out\[10\] net1876 _01003_ VPWR VGND sg13g2_mux2_1
XFILLER_46_736 VPWR VGND sg13g2_decap_8
XFILLER_18_438 VPWR VGND sg13g2_decap_4
XFILLER_61_717 VPWR VGND sg13g2_fill_1
X_14620_ _00421_ VGND VPWR _01152_ fp16_sum_pipe.exp_mant_logic0.a\[15\] clknet_leaf_124_clk
+ sg13g2_dfrbpq_2
X_11832_ VGND VPWR _05638_ _05639_ _05731_ _05489_ sg13g2_a21oi_1
X_14551_ _00352_ VGND VPWR _01087_ acc_sum.op_sign_logic0.mantisa_a\[3\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_61_739 VPWR VGND sg13g2_fill_1
XFILLER_60_238 VPWR VGND sg13g2_decap_8
XFILLER_45_279 VPWR VGND sg13g2_decap_8
XFILLER_14_611 VPWR VGND sg13g2_decap_8
XFILLER_14_622 VPWR VGND sg13g2_fill_2
XFILLER_26_84 VPWR VGND sg13g2_decap_8
XFILLER_42_964 VPWR VGND sg13g2_decap_8
XFILLER_41_441 VPWR VGND sg13g2_decap_8
XFILLER_13_132 VPWR VGND sg13g2_decap_8
X_11763_ _05662_ _05666_ _05667_ VPWR VGND sg13g2_nor2_1
X_13502_ VPWR _00053_ net90 VGND sg13g2_inv_1
XFILLER_42_997 VPWR VGND sg13g2_decap_4
X_14482_ _00283_ VGND VPWR _01020_ add_result\[7\] clknet_leaf_98_clk sg13g2_dfrbpq_1
X_10714_ _04727_ _04726_ _04695_ VPWR VGND sg13g2_nand2_1
X_11694_ _05598_ _05596_ VPWR VGND sg13g2_inv_2
X_13433_ _07095_ VPWR _00787_ VGND _07018_ net1720 sg13g2_o21ai_1
XFILLER_9_147 VPWR VGND sg13g2_decap_4
X_10645_ _04655_ _04657_ _04658_ VPWR VGND sg13g2_nor2b_2
XFILLER_127_513 VPWR VGND sg13g2_decap_8
XFILLER_61_9 VPWR VGND sg13g2_fill_1
X_12315_ _06161_ net1860 net1865 VPWR VGND sg13g2_nand2_1
X_10576_ _04601_ acc_sub.x2\[11\] net1924 VPWR VGND sg13g2_nand2_1
XFILLER_6_843 VPWR VGND sg13g2_decap_8
XFILLER_114_207 VPWR VGND sg13g2_decap_8
XFILLER_108_771 VPWR VGND sg13g2_decap_8
X_13295_ acc\[4\] net1678 _07009_ VPWR VGND sg13g2_nor2_1
XFILLER_108_782 VPWR VGND sg13g2_fill_2
X_12246_ _06090_ _06091_ _06092_ VPWR VGND sg13g2_nor2_2
XFILLER_5_386 VPWR VGND sg13g2_decap_8
X_12177_ VGND VPWR _06007_ _05983_ _06023_ _06022_ sg13g2_a21oi_1
XFILLER_123_785 VPWR VGND sg13g2_decap_8
XFILLER_122_273 VPWR VGND sg13g2_decap_8
XFILLER_111_936 VPWR VGND sg13g2_decap_8
XFILLER_95_113 VPWR VGND sg13g2_fill_1
X_11128_ _05098_ _05006_ _05097_ VPWR VGND sg13g2_xnor2_1
XFILLER_3_77 VPWR VGND sg13g2_decap_8
XFILLER_95_168 VPWR VGND sg13g2_fill_1
XFILLER_77_883 VPWR VGND sg13g2_fill_1
X_11059_ VPWR _05037_ _05003_ VGND sg13g2_inv_1
XFILLER_36_202 VPWR VGND sg13g2_fill_1
XFILLER_36_235 VPWR VGND sg13g2_decap_8
X_14818_ _00619_ VGND VPWR _01342_ acc_sum.add_renorm0.mantisa\[7\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_64_555 VPWR VGND sg13g2_fill_2
XFILLER_58_1008 VPWR VGND sg13g2_decap_4
XFILLER_91_385 VPWR VGND sg13g2_decap_8
XFILLER_18_983 VPWR VGND sg13g2_decap_8
X_14749_ _00550_ VGND VPWR _01277_ fp16_res_pipe.seg_reg1.q\[20\] clknet_leaf_130_clk
+ sg13g2_dfrbpq_1
XFILLER_33_953 VPWR VGND sg13g2_decap_8
X_08270_ _02519_ _02408_ _02472_ VPWR VGND sg13g2_nand2_1
XFILLER_20_625 VPWR VGND sg13g2_decap_8
XFILLER_32_463 VPWR VGND sg13g2_fill_1
XFILLER_20_647 VPWR VGND sg13g2_decap_8
X_07152_ acc_sub.op_sign_logic0.mantisa_b\[6\] _01523_ _01524_ VPWR VGND sg13g2_nor2_1
XFILLER_73_0 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_8_clk clknet_5_4__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
XFILLER_114_730 VPWR VGND sg13g2_fill_1
XFILLER_99_430 VPWR VGND sg13g2_decap_8
XFILLER_114_741 VPWR VGND sg13g2_decap_8
Xfanout104 net107 net104 VPWR VGND sg13g2_buf_1
XFILLER_87_603 VPWR VGND sg13g2_fill_1
XFILLER_99_485 VPWR VGND sg13g2_fill_1
Xfanout137 net138 net137 VPWR VGND sg13g2_buf_2
Xfanout126 net127 net126 VPWR VGND sg13g2_buf_1
XFILLER_87_614 VPWR VGND sg13g2_decap_8
Xfanout115 net116 net115 VPWR VGND sg13g2_buf_1
XFILLER_113_295 VPWR VGND sg13g2_decap_8
XFILLER_102_958 VPWR VGND sg13g2_decap_8
XFILLER_86_146 VPWR VGND sg13g2_fill_2
X_07985_ _02255_ VPWR _01387_ VGND _02205_ _02248_ sg13g2_o21ai_1
X_09724_ _03840_ _02930_ _03839_ VPWR VGND sg13g2_xnor2_1
XFILLER_68_883 VPWR VGND sg13g2_decap_8
XFILLER_55_500 VPWR VGND sg13g2_decap_8
X_09655_ _03732_ _03771_ _03730_ _03772_ VPWR VGND sg13g2_nand3_1
XFILLER_67_371 VPWR VGND sg13g2_fill_1
X_08606_ _02829_ _02828_ net1739 VPWR VGND sg13g2_nand2_1
XFILLER_82_341 VPWR VGND sg13g2_decap_8
XFILLER_27_246 VPWR VGND sg13g2_decap_4
X_09586_ _03702_ VPWR _03703_ VGND _02806_ acc_sum.add_renorm0.mantisa\[4\] sg13g2_o21ai_1
XFILLER_83_897 VPWR VGND sg13g2_decap_8
X_08537_ VPWR _02761_ acc_sum.op_sign_logic0.mantisa_b\[0\] VGND sg13g2_inv_1
XFILLER_24_953 VPWR VGND sg13g2_decap_8
X_08468_ _02699_ VPWR _02700_ VGND fpdiv.divider0.remainder_reg\[9\] net1647 sg13g2_o21ai_1
XFILLER_23_474 VPWR VGND sg13g2_decap_8
X_07419_ _01754_ VPWR _01452_ VGND net1890 _01753_ sg13g2_o21ai_1
XFILLER_50_293 VPWR VGND sg13g2_fill_2
XFILLER_23_485 VPWR VGND sg13g2_fill_1
X_08399_ _02636_ _02589_ state\[1\] VPWR VGND sg13g2_nand2_1
X_10430_ _04479_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[2\] fp16_sum_pipe.op_sign_logic0.mantisa_b\[2\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_109_546 VPWR VGND sg13g2_fill_2
XFILLER_12_42 VPWR VGND sg13g2_decap_8
XFILLER_109_579 VPWR VGND sg13g2_decap_4
X_10361_ VPWR _04411_ _04410_ VGND sg13g2_inv_1
X_13080_ VGND VPWR _06811_ _06759_ _06845_ _06835_ sg13g2_a21oi_1
X_12100_ _05898_ _05905_ _05942_ _05946_ VPWR VGND sg13g2_nand3_1
X_10292_ _04360_ fp16_res_pipe.exp_mant_logic0.b\[4\] _04210_ _04224_ net1830 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_88_68 VPWR VGND sg13g2_fill_1
XFILLER_88_57 VPWR VGND sg13g2_fill_1
X_12031_ _05878_ fpmul.reg_a_out\[7\] fpmul.reg_b_out\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_3_868 VPWR VGND sg13g2_decap_8
XFILLER_120_711 VPWR VGND sg13g2_decap_8
XFILLER_78_625 VPWR VGND sg13g2_fill_2
XFILLER_2_367 VPWR VGND sg13g2_decap_8
XFILLER_120_799 VPWR VGND sg13g2_decap_8
X_13982_ VPWR _00533_ net13 VGND sg13g2_inv_1
XFILLER_86_680 VPWR VGND sg13g2_decap_8
X_12933_ acc\[3\] net1907 _03983_ _06706_ VPWR VGND sg13g2_nand3_1
XFILLER_46_533 VPWR VGND sg13g2_fill_1
XFILLER_46_522 VPWR VGND sg13g2_decap_8
XFILLER_19_725 VPWR VGND sg13g2_decap_4
XFILLER_74_864 VPWR VGND sg13g2_fill_1
X_12864_ _06643_ _06639_ _06642_ _06496_ net1943 VPWR VGND sg13g2_a22oi_1
XFILLER_15_931 VPWR VGND sg13g2_decap_8
XFILLER_33_205 VPWR VGND sg13g2_decap_4
XFILLER_61_547 VPWR VGND sg13g2_decap_4
X_14603_ _00404_ VGND VPWR _01135_ fp16_res_pipe.y\[14\] clknet_leaf_129_clk sg13g2_dfrbpq_1
X_11815_ _05716_ _05706_ _05715_ VPWR VGND sg13g2_nand2_1
X_14534_ _00335_ VGND VPWR _01070_ fpdiv.div_out\[9\] clknet_leaf_77_clk sg13g2_dfrbpq_1
X_11746_ _05650_ _05631_ _05649_ VPWR VGND sg13g2_nand2_1
XFILLER_53_82 VPWR VGND sg13g2_decap_8
XFILLER_30_934 VPWR VGND sg13g2_decap_8
X_14465_ _00266_ VGND VPWR _01004_ fpmul.seg_reg0.q\[50\] clknet_leaf_96_clk sg13g2_dfrbpq_1
X_11677_ _05581_ _04581_ _05580_ VPWR VGND sg13g2_xnor2_1
X_14396_ _00197_ VGND VPWR _00935_ div_result\[9\] clknet_leaf_89_clk sg13g2_dfrbpq_1
X_13416_ _07087_ net1722 instr\[9\] VPWR VGND sg13g2_nand2_1
X_10628_ _04641_ fp16_res_pipe.add_renorm0.mantisa\[3\] fp16_res_pipe.add_renorm0.mantisa\[2\]
+ VPWR VGND sg13g2_nand2_1
XFILLER_127_343 VPWR VGND sg13g2_decap_8
Xplace1818 net1816 net1818 VPWR VGND sg13g2_buf_2
Xplace1807 acc_sum.add_renorm0.mantisa\[11\] net1807 VPWR VGND sg13g2_buf_2
X_13347_ _07047_ VPWR _00825_ VGND _07046_ _07027_ sg13g2_o21ai_1
X_10559_ VPWR _04591_ fp16_sum_pipe.add_renorm0.exp\[2\] VGND sg13g2_inv_1
X_13278_ acc\[8\] _06995_ net1678 _00842_ VPWR VGND sg13g2_mux2_1
XFILLER_5_161 VPWR VGND sg13g2_decap_8
Xplace1829 fp16_res_pipe.exp_mant_logic0.b\[6\] net1829 VPWR VGND sg13g2_buf_2
X_12229_ _06075_ _06072_ _06074_ VPWR VGND sg13g2_xnor2_1
XFILLER_123_560 VPWR VGND sg13g2_decap_8
XFILLER_111_722 VPWR VGND sg13g2_decap_8
XFILLER_97_956 VPWR VGND sg13g2_decap_8
X_07770_ _02072_ net1795 net1669 acc_sub.op_sign_logic0.mantisa_b\[8\] net1781 VPWR
+ VGND sg13g2_a22oi_1
XFILLER_84_628 VPWR VGND sg13g2_decap_8
XFILLER_68_168 VPWR VGND sg13g2_decap_8
XFILLER_96_499 VPWR VGND sg13g2_decap_8
XFILLER_84_639 VPWR VGND sg13g2_fill_1
XFILLER_83_138 VPWR VGND sg13g2_decap_8
XFILLER_77_680 VPWR VGND sg13g2_fill_2
X_09440_ _03579_ net1834 fp16_res_pipe.seg_reg0.q\[27\] VPWR VGND sg13g2_nand2_1
XFILLER_92_694 VPWR VGND sg13g2_fill_1
XFILLER_64_363 VPWR VGND sg13g2_decap_8
XFILLER_91_193 VPWR VGND sg13g2_decap_8
X_09371_ _03520_ VPWR _01273_ VGND fp16_res_pipe.reg2en.q\[0\] _03512_ sg13g2_o21ai_1
X_08322_ VPWR _02567_ state\[0\] VGND sg13g2_inv_1
X_08253_ _02504_ net1638 _02503_ VPWR VGND sg13g2_nand2_1
XFILLER_21_945 VPWR VGND sg13g2_decap_8
XFILLER_32_260 VPWR VGND sg13g2_decap_8
XFILLER_119_800 VPWR VGND sg13g2_decap_8
X_07204_ VGND VPWR _01521_ _01524_ _01576_ _01518_ sg13g2_a21oi_1
X_08184_ _02438_ _02441_ _02437_ _02442_ VPWR VGND sg13g2_nand3_1
XFILLER_119_877 VPWR VGND sg13g2_decap_8
X_07135_ _01504_ _01506_ _01507_ VPWR VGND sg13g2_nor2_2
XFILLER_121_519 VPWR VGND sg13g2_fill_1
XFILLER_102_722 VPWR VGND sg13g2_decap_8
XFILLER_114_593 VPWR VGND sg13g2_decap_8
XFILLER_88_967 VPWR VGND sg13g2_decap_8
XFILLER_58_49 VPWR VGND sg13g2_decap_4
XFILLER_0_849 VPWR VGND sg13g2_decap_8
XFILLER_102_777 VPWR VGND sg13g2_decap_4
XFILLER_75_628 VPWR VGND sg13g2_fill_2
XFILLER_74_105 VPWR VGND sg13g2_fill_1
X_07968_ VGND VPWR _02241_ _02186_ _02242_ _02179_ sg13g2_a21oi_1
X_09707_ _03823_ _03819_ _03822_ VPWR VGND sg13g2_nand2_1
XFILLER_87_499 VPWR VGND sg13g2_decap_8
XFILLER_28_533 VPWR VGND sg13g2_fill_1
XFILLER_114_77 VPWR VGND sg13g2_decap_8
X_07899_ _02176_ VPWR _01394_ VGND net1892 _02130_ sg13g2_o21ai_1
XFILLER_83_661 VPWR VGND sg13g2_fill_2
XFILLER_74_37 VPWR VGND sg13g2_decap_8
XFILLER_16_706 VPWR VGND sg13g2_decap_8
XFILLER_28_555 VPWR VGND sg13g2_decap_4
X_09638_ _03753_ _03754_ _03752_ _03755_ VPWR VGND sg13g2_nand3_1
XFILLER_70_300 VPWR VGND sg13g2_decap_4
X_09569_ _03686_ _03635_ _03666_ _03641_ _03630_ VPWR VGND sg13g2_a22oi_1
XFILLER_15_227 VPWR VGND sg13g2_decap_4
X_12580_ _06389_ _06392_ _06396_ VPWR VGND sg13g2_xor2_1
XFILLER_70_377 VPWR VGND sg13g2_decap_4
X_11600_ _05504_ VPWR _05505_ VGND _05502_ _05503_ sg13g2_o21ai_1
XFILLER_30_219 VPWR VGND sg13g2_decap_8
XFILLER_90_47 VPWR VGND sg13g2_fill_2
XFILLER_11_433 VPWR VGND sg13g2_decap_8
X_11531_ VPWR _05436_ fp16_sum_pipe.add_renorm0.mantisa\[8\] VGND sg13g2_inv_1
XFILLER_23_260 VPWR VGND sg13g2_decap_8
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_12_967 VPWR VGND sg13g2_decap_8
XFILLER_23_63 VPWR VGND sg13g2_decap_8
XFILLER_109_332 VPWR VGND sg13g2_decap_4
X_11462_ _05384_ acc_sub.x2\[0\] net1947 VPWR VGND sg13g2_nand2_1
X_14250_ _00051_ VGND VPWR _00801_ instr\[15\] clknet_leaf_15_clk sg13g2_dfrbpq_1
XFILLER_11_488 VPWR VGND sg13g2_decap_8
X_14181_ VPWR _00732_ net139 VGND sg13g2_inv_1
XFILLER_99_23 VPWR VGND sg13g2_fill_1
X_11393_ _05340_ VPWR _01071_ VGND _05339_ net1706 sg13g2_o21ai_1
X_13201_ VPWR _06935_ sipo.shift_reg\[4\] VGND sg13g2_inv_1
X_10413_ VGND VPWR _04460_ _02177_ _04463_ _04462_ sg13g2_a21oi_1
XFILLER_125_858 VPWR VGND sg13g2_decap_8
XFILLER_109_387 VPWR VGND sg13g2_fill_2
XFILLER_99_67 VPWR VGND sg13g2_decap_8
X_13132_ VGND VPWR _06882_ _06570_ _06884_ piso.tx_bit_counter\[3\] sg13g2_a21oi_1
X_10344_ fp16_sum_pipe.op_sign_logic0.mantisa_b\[9\] _04393_ _04394_ VPWR VGND sg13g2_nor2_1
XFILLER_3_0 VPWR VGND sg13g2_decap_8
X_13063_ _05795_ _05797_ _05793_ _06831_ VPWR VGND _05799_ sg13g2_nand4_1
X_10275_ _04342_ _04344_ _04345_ VPWR VGND sg13g2_nor2_1
X_12014_ _05865_ VPWR _00975_ VGND net1877 _05863_ sg13g2_o21ai_1
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_120_574 VPWR VGND sg13g2_fill_1
XFILLER_120_552 VPWR VGND sg13g2_fill_1
XFILLER_94_926 VPWR VGND sg13g2_decap_8
XFILLER_66_628 VPWR VGND sg13g2_fill_2
XFILLER_66_617 VPWR VGND sg13g2_decap_8
XFILLER_65_138 VPWR VGND sg13g2_decap_8
XFILLER_19_511 VPWR VGND sg13g2_decap_8
X_13965_ VPWR _00516_ net7 VGND sg13g2_inv_1
XFILLER_80_119 VPWR VGND sg13g2_decap_4
X_12916_ _06691_ _06690_ net1733 VPWR VGND sg13g2_nand2_1
XFILLER_62_834 VPWR VGND sg13g2_decap_4
XFILLER_47_886 VPWR VGND sg13g2_fill_2
XFILLER_46_374 VPWR VGND sg13g2_decap_8
X_13896_ VPWR _00447_ net17 VGND sg13g2_inv_1
XFILLER_0_56 VPWR VGND sg13g2_decap_8
X_12847_ VPWR _06627_ div_result\[10\] VGND sg13g2_inv_1
XFILLER_61_322 VPWR VGND sg13g2_decap_8
XFILLER_61_377 VPWR VGND sg13g2_fill_2
XFILLER_61_355 VPWR VGND sg13g2_fill_2
XFILLER_9_21 VPWR VGND sg13g2_decap_8
X_12778_ _06562_ VPWR _06563_ VGND net1958 _06551_ sg13g2_o21ai_1
X_14517_ _00318_ VGND VPWR _01053_ fpdiv.reg_a_out\[8\] clknet_leaf_91_clk sg13g2_dfrbpq_2
X_11729_ _05633_ _05632_ _05596_ VPWR VGND sg13g2_nand2_1
X_14448_ _00249_ VGND VPWR _00987_ fpmul.seg_reg0.q\[33\] clknet_leaf_97_clk sg13g2_dfrbpq_1
XFILLER_9_98 VPWR VGND sg13g2_decap_8
XFILLER_127_140 VPWR VGND sg13g2_decap_8
XFILLER_116_814 VPWR VGND sg13g2_decap_8
X_14379_ _00180_ VGND VPWR _00920_ fpmul.reg_b_out\[10\] clknet_leaf_124_clk sg13g2_dfrbpq_2
XFILLER_7_993 VPWR VGND sg13g2_decap_8
XFILLER_6_481 VPWR VGND sg13g2_decap_8
XFILLER_89_709 VPWR VGND sg13g2_fill_1
Xplace1659 _02338_ net1659 VPWR VGND sg13g2_buf_1
Xplace1648 _02345_ net1648 VPWR VGND sg13g2_buf_1
Xplace1637 _04150_ net1637 VPWR VGND sg13g2_buf_2
X_08940_ _03127_ _03009_ _03004_ VPWR VGND sg13g2_nand2_1
XFILLER_69_400 VPWR VGND sg13g2_decap_4
X_08871_ _03031_ _03057_ _03058_ VPWR VGND sg13g2_nor2_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
XFILLER_111_552 VPWR VGND sg13g2_decap_8
X_07822_ _02114_ _02118_ _02119_ VPWR VGND sg13g2_nor2_1
XFILLER_84_403 VPWR VGND sg13g2_fill_2
XFILLER_96_285 VPWR VGND sg13g2_decap_4
XFILLER_84_436 VPWR VGND sg13g2_decap_8
XFILLER_57_639 VPWR VGND sg13g2_decap_8
X_07753_ acc_sub.exp_mant_logic0.b\[2\] acc_sub.exp_mant_logic0.b\[1\] acc_sub.exp_mant_logic0.b\[0\]
+ _02057_ VPWR VGND sg13g2_nor3_1
X_07684_ VGND VPWR net1793 _01935_ _01993_ _01992_ sg13g2_a21oi_1
XFILLER_65_694 VPWR VGND sg13g2_decap_4
XFILLER_65_683 VPWR VGND sg13g2_decap_8
XFILLER_38_897 VPWR VGND sg13g2_decap_8
XFILLER_80_631 VPWR VGND sg13g2_decap_4
XFILLER_53_856 VPWR VGND sg13g2_fill_1
X_09423_ _03566_ _03459_ _03443_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_558 VPWR VGND sg13g2_decap_8
XFILLER_53_878 VPWR VGND sg13g2_fill_1
X_09354_ _03505_ net1770 fp16_res_pipe.add_renorm0.mantisa\[9\] VPWR VGND sg13g2_nand2_1
X_08305_ _01363_ _02550_ _02551_ VPWR VGND sg13g2_nand2_1
XFILLER_100_68 VPWR VGND sg13g2_decap_8
X_09285_ VPWR VGND _03438_ _03373_ _03433_ _03371_ _03439_ _03377_ sg13g2_a221oi_1
X_08236_ _02489_ net1638 _02488_ VPWR VGND sg13g2_nand2_1
XFILLER_118_140 VPWR VGND sg13g2_decap_8
XFILLER_107_803 VPWR VGND sg13g2_fill_1
X_08167_ _02336_ _02327_ _02426_ VPWR VGND sg13g2_nor2_1
XFILLER_114_7 VPWR VGND sg13g2_decap_8
XFILLER_106_324 VPWR VGND sg13g2_fill_2
XFILLER_109_77 VPWR VGND sg13g2_fill_2
XFILLER_107_858 VPWR VGND sg13g2_decap_8
X_08098_ _01381_ _02361_ _02362_ VPWR VGND sg13g2_nand2_1
XFILLER_106_368 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_fill_1
XFILLER_0_613 VPWR VGND sg13g2_decap_8
XFILLER_125_21 VPWR VGND sg13g2_decap_8
XFILLER_87_230 VPWR VGND sg13g2_decap_8
X_10060_ _04148_ _04140_ _04147_ VPWR VGND sg13g2_nand2_1
XFILLER_88_775 VPWR VGND sg13g2_decap_8
XFILLER_125_98 VPWR VGND sg13g2_decap_8
XFILLER_48_639 VPWR VGND sg13g2_decap_4
XFILLER_48_628 VPWR VGND sg13g2_fill_2
XFILLER_56_650 VPWR VGND sg13g2_decap_8
XFILLER_47_138 VPWR VGND sg13g2_fill_2
X_13750_ VPWR _00301_ net115 VGND sg13g2_inv_1
XFILLER_56_683 VPWR VGND sg13g2_fill_1
XFILLER_43_300 VPWR VGND sg13g2_fill_2
X_10962_ _04967_ _04772_ fp16_res_pipe.y\[7\] VPWR VGND sg13g2_nand2_1
XFILLER_18_63 VPWR VGND sg13g2_decap_8
X_12701_ _06509_ VPWR _00933_ VGND _06502_ net1741 sg13g2_o21ai_1
X_13681_ VPWR _00232_ net69 VGND sg13g2_inv_1
XFILLER_43_355 VPWR VGND sg13g2_fill_2
X_10893_ _04796_ _04850_ _04903_ VPWR VGND sg13g2_nor2_1
X_12632_ _06448_ _06443_ _06447_ VPWR VGND sg13g2_nand2_1
X_12563_ _06379_ _05389_ fpdiv.reg_a_out\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_34_84 VPWR VGND sg13g2_decap_8
XFILLER_11_230 VPWR VGND sg13g2_decap_4
XFILLER_12_753 VPWR VGND sg13g2_decap_8
X_14302_ _00103_ VGND VPWR _00846_ acc\[12\] clknet_leaf_49_clk sg13g2_dfrbpq_2
X_12494_ VGND VPWR _06328_ net1871 _00959_ _06329_ sg13g2_a21oi_1
XFILLER_8_746 VPWR VGND sg13g2_decap_8
XFILLER_11_252 VPWR VGND sg13g2_decap_8
X_11514_ _05419_ fp16_sum_pipe.add_renorm0.mantisa\[6\] VPWR VGND sg13g2_inv_2
X_11445_ _05373_ acc_sub.x2\[6\] net1946 VPWR VGND sg13g2_nand2_1
X_14233_ _00034_ VGND VPWR _00784_ sipo.shift_reg\[14\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_14164_ VPWR _00715_ net102 VGND sg13g2_inv_1
X_11376_ _05325_ _05326_ _05327_ VPWR VGND sg13g2_nor2b_1
XFILLER_4_930 VPWR VGND sg13g2_decap_8
XFILLER_125_688 VPWR VGND sg13g2_fill_2
XFILLER_124_154 VPWR VGND sg13g2_decap_8
X_13115_ net1700 _06871_ _06802_ _06872_ VPWR VGND sg13g2_nand3_1
X_14095_ VPWR _00646_ net40 VGND sg13g2_inv_1
XFILLER_3_462 VPWR VGND sg13g2_decap_8
X_10327_ _04381_ net1921 fp16_res_pipe.x2\[2\] VPWR VGND sg13g2_nand2_1
X_13046_ _06757_ _06813_ _06814_ VPWR VGND sg13g2_nor2_1
X_10258_ _04329_ fp16_res_pipe.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_inv_2
XFILLER_121_861 VPWR VGND sg13g2_decap_8
XFILLER_67_915 VPWR VGND sg13g2_decap_8
XFILLER_93_200 VPWR VGND sg13g2_decap_8
XFILLER_39_639 VPWR VGND sg13g2_fill_1
XFILLER_39_628 VPWR VGND sg13g2_fill_2
XFILLER_38_105 VPWR VGND sg13g2_decap_8
X_10189_ fp16_res_pipe.exp_mant_logic0.b\[2\] fp16_res_pipe.exp_mant_logic0.b\[1\]
+ fp16_res_pipe.exp_mant_logic0.b\[0\] _04267_ VPWR VGND sg13g2_nor3_1
XFILLER_93_255 VPWR VGND sg13g2_decap_8
XFILLER_66_458 VPWR VGND sg13g2_decap_8
XFILLER_47_650 VPWR VGND sg13g2_fill_1
X_13948_ VPWR _00499_ net97 VGND sg13g2_inv_1
XFILLER_53_108 VPWR VGND sg13g2_decap_4
XFILLER_46_160 VPWR VGND sg13g2_decap_8
XFILLER_35_812 VPWR VGND sg13g2_decap_8
XFILLER_34_311 VPWR VGND sg13g2_decap_8
XFILLER_19_396 VPWR VGND sg13g2_fill_2
XFILLER_90_995 VPWR VGND sg13g2_decap_8
XFILLER_62_686 VPWR VGND sg13g2_decap_8
X_13879_ VPWR _00430_ net48 VGND sg13g2_inv_1
XFILLER_50_848 VPWR VGND sg13g2_fill_2
XFILLER_22_539 VPWR VGND sg13g2_fill_2
X_09070_ _03255_ _03247_ _03254_ VPWR VGND sg13g2_nand2_1
X_08021_ _02189_ _02286_ _02187_ _02287_ VPWR VGND sg13g2_a21o_1
Xfanout6 net15 net6 VPWR VGND sg13g2_buf_1
XFILLER_115_154 VPWR VGND sg13g2_decap_8
XFILLER_103_305 VPWR VGND sg13g2_decap_8
X_09972_ _04064_ net1765 fp16_res_pipe.seg_reg0.q\[24\] VPWR VGND sg13g2_nand2_1
X_08923_ _03110_ _03042_ _03021_ VPWR VGND sg13g2_nand2_1
X_08854_ _03040_ VPWR _03041_ VGND net1789 _02982_ sg13g2_o21ai_1
XFILLER_112_894 VPWR VGND sg13g2_decap_8
XFILLER_111_360 VPWR VGND sg13g2_decap_8
XFILLER_97_583 VPWR VGND sg13g2_decap_4
XFILLER_69_296 VPWR VGND sg13g2_decap_8
X_07805_ _02103_ net1650 net1795 VPWR VGND sg13g2_nand2_1
XFILLER_85_767 VPWR VGND sg13g2_decap_8
XFILLER_73_918 VPWR VGND sg13g2_decap_8
XFILLER_45_609 VPWR VGND sg13g2_fill_2
X_07736_ _01422_ _02040_ _02041_ VPWR VGND sg13g2_nand2_1
XFILLER_55_28 VPWR VGND sg13g2_decap_8
XFILLER_44_119 VPWR VGND sg13g2_decap_8
XFILLER_26_856 VPWR VGND sg13g2_decap_8
XFILLER_111_56 VPWR VGND sg13g2_decap_8
X_07667_ _01977_ _01975_ VPWR VGND sg13g2_inv_2
XFILLER_52_130 VPWR VGND sg13g2_decap_8
X_07598_ _01911_ VPWR _01912_ VGND _01827_ net1686 sg13g2_o21ai_1
X_09406_ _03551_ net1675 _03490_ VPWR VGND sg13g2_nand2_1
XFILLER_25_399 VPWR VGND sg13g2_fill_2
X_09337_ VPWR _03489_ _03488_ VGND sg13g2_inv_1
X_09268_ fp16_res_pipe.op_sign_logic0.mantisa_a\[4\] _03421_ _03422_ VPWR VGND sg13g2_nor2_1
XFILLER_21_561 VPWR VGND sg13g2_fill_1
X_08219_ _02474_ _02472_ net1645 net1691 fp16_sum_pipe.exp_mant_logic0.b\[6\] VPWR
+ VGND sg13g2_a22oi_1
XFILLER_107_600 VPWR VGND sg13g2_decap_4
X_09199_ _03356_ acc_sub.x2\[1\] net1905 VPWR VGND sg13g2_nand2_1
XFILLER_106_121 VPWR VGND sg13g2_fill_1
X_11230_ _05072_ _05194_ _05195_ VPWR VGND sg13g2_nor2_1
XFILLER_20_42 VPWR VGND sg13g2_decap_8
XFILLER_106_165 VPWR VGND sg13g2_decap_8
X_11161_ VPWR _05130_ _05106_ VGND sg13g2_inv_1
XFILLER_20_86 VPWR VGND sg13g2_fill_2
XFILLER_0_421 VPWR VGND sg13g2_decap_8
X_10112_ _04143_ _04131_ _04195_ VPWR VGND sg13g2_nor2_2
XFILLER_121_168 VPWR VGND sg13g2_decap_8
X_11092_ _05065_ _05052_ acc_sum.exp_mant_logic0.a\[8\] VPWR VGND sg13g2_nand2_1
XFILLER_1_955 VPWR VGND sg13g2_decap_8
X_14920_ _00721_ VGND VPWR _01440_ acc_sub.op_sign_logic0.add_sub clknet_leaf_62_clk
+ sg13g2_dfrbpq_2
XFILLER_88_572 VPWR VGND sg13g2_decap_4
X_10043_ _04097_ _04103_ _04131_ VPWR VGND _04090_ sg13g2_nand3b_1
XFILLER_0_498 VPWR VGND sg13g2_decap_8
X_14851_ _00652_ VGND VPWR _01375_ fp16_sum_pipe.op_sign_logic0.mantisa_a\[2\] clknet_leaf_114_clk
+ sg13g2_dfrbpq_2
XFILLER_91_737 VPWR VGND sg13g2_decap_4
XFILLER_91_726 VPWR VGND sg13g2_fill_1
XFILLER_90_203 VPWR VGND sg13g2_decap_4
X_13802_ VPWR _00353_ net73 VGND sg13g2_inv_1
XFILLER_63_428 VPWR VGND sg13g2_decap_4
XFILLER_63_417 VPWR VGND sg13g2_fill_2
XFILLER_57_981 VPWR VGND sg13g2_fill_1
XFILLER_35_119 VPWR VGND sg13g2_decap_8
XFILLER_17_812 VPWR VGND sg13g2_fill_2
X_14782_ _00583_ VGND VPWR _01306_ acc_sub.y\[11\] clknet_leaf_38_clk sg13g2_dfrbpq_1
X_11994_ _05848_ _05831_ _05829_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_856 VPWR VGND sg13g2_decap_8
XFILLER_72_984 VPWR VGND sg13g2_decap_8
X_13733_ VPWR _00284_ net63 VGND sg13g2_inv_1
XFILLER_44_675 VPWR VGND sg13g2_decap_8
XFILLER_44_653 VPWR VGND sg13g2_fill_1
XFILLER_16_366 VPWR VGND sg13g2_decap_4
X_10945_ _04951_ _04843_ _04842_ VPWR VGND sg13g2_nand2_1
XFILLER_32_804 VPWR VGND sg13g2_decap_8
XFILLER_72_995 VPWR VGND sg13g2_fill_1
X_13664_ VPWR _00215_ net57 VGND sg13g2_inv_1
XFILLER_16_399 VPWR VGND sg13g2_fill_2
X_10876_ _04887_ _04826_ _04849_ VPWR VGND sg13g2_nand2_1
XFILLER_32_848 VPWR VGND sg13g2_decap_8
XFILLER_32_859 VPWR VGND sg13g2_fill_1
X_12615_ _06431_ _06425_ _06429_ _06430_ VPWR VGND sg13g2_and3_1
X_13595_ VPWR _00146_ net110 VGND sg13g2_inv_1
XFILLER_12_561 VPWR VGND sg13g2_decap_8
XFILLER_12_572 VPWR VGND sg13g2_fill_1
X_12546_ _06363_ _06361_ _06362_ VPWR VGND sg13g2_nand2_1
XFILLER_77_7 VPWR VGND sg13g2_fill_1
XFILLER_12_583 VPWR VGND sg13g2_fill_1
X_12477_ _06316_ _06149_ _06317_ VPWR VGND sg13g2_xor2_1
XFILLER_8_587 VPWR VGND sg13g2_fill_2
XFILLER_126_953 VPWR VGND sg13g2_decap_8
X_14216_ VPWR _00767_ net132 VGND sg13g2_inv_1
X_11428_ _05362_ acc_sub.x2\[12\] net1938 VPWR VGND sg13g2_nand2_1
XFILLER_125_463 VPWR VGND sg13g2_fill_2
X_14147_ VPWR _00698_ net134 VGND sg13g2_inv_1
XFILLER_113_614 VPWR VGND sg13g2_decap_4
X_11359_ _05311_ _05146_ acc_sum.exp_mant_logic0.b\[3\] VPWR VGND sg13g2_nand2_1
XFILLER_6_77 VPWR VGND sg13g2_decap_8
XFILLER_99_859 VPWR VGND sg13g2_fill_2
X_14078_ VPWR _00629_ net138 VGND sg13g2_inv_1
XFILLER_94_520 VPWR VGND sg13g2_decap_8
X_13029_ _06797_ net1853 fpmul.seg_reg0.q\[6\] VPWR VGND sg13g2_nand2_1
XFILLER_39_425 VPWR VGND sg13g2_decap_8
XFILLER_39_414 VPWR VGND sg13g2_decap_8
XFILLER_6_1004 VPWR VGND sg13g2_decap_8
XFILLER_66_244 VPWR VGND sg13g2_decap_8
XFILLER_66_222 VPWR VGND sg13g2_fill_1
XFILLER_39_447 VPWR VGND sg13g2_decap_8
XFILLER_39_436 VPWR VGND sg13g2_fill_1
XFILLER_27_609 VPWR VGND sg13g2_decap_4
X_08570_ VPWR _02794_ _02793_ VGND sg13g2_inv_1
XFILLER_82_726 VPWR VGND sg13g2_decap_8
XFILLER_26_108 VPWR VGND sg13g2_decap_8
X_07452_ net1796 acc_sub.op_sign_logic0.s_b _01777_ VPWR VGND sg13g2_nor2_1
XFILLER_63_995 VPWR VGND sg13g2_decap_4
X_07383_ _01730_ VPWR _01464_ VGND net1886 _01729_ sg13g2_o21ai_1
XFILLER_50_656 VPWR VGND sg13g2_decap_8
X_09122_ net1786 VPWR _03303_ VGND _03229_ _03302_ sg13g2_o21ai_1
X_09053_ VGND VPWR _03151_ net1791 _03239_ _03238_ sg13g2_a21oi_1
XFILLER_117_942 VPWR VGND sg13g2_decap_8
X_08004_ _02268_ _02269_ _02267_ _02271_ VPWR VGND _02270_ sg13g2_nand4_1
XFILLER_89_303 VPWR VGND sg13g2_fill_2
XFILLER_106_23 VPWR VGND sg13g2_fill_2
X_09955_ _04050_ _04047_ _04029_ VPWR VGND sg13g2_nand2_2
X_08906_ _03092_ _02996_ _03083_ _03093_ VPWR VGND sg13g2_nor3_1
XFILLER_57_200 VPWR VGND sg13g2_fill_2
X_09886_ VPWR _03985_ fp16_res_pipe.exp_mant_logic0.b\[15\] VGND sg13g2_inv_1
X_08837_ VPWR _03024_ net1788 VGND sg13g2_inv_1
XFILLER_100_853 VPWR VGND sg13g2_fill_1
XFILLER_100_831 VPWR VGND sg13g2_fill_1
XFILLER_66_49 VPWR VGND sg13g2_fill_2
XFILLER_58_756 VPWR VGND sg13g2_decap_8
XFILLER_73_726 VPWR VGND sg13g2_fill_1
XFILLER_58_789 VPWR VGND sg13g2_decap_8
XFILLER_58_778 VPWR VGND sg13g2_fill_1
XFILLER_39_970 VPWR VGND sg13g2_decap_8
X_08768_ _02958_ VPWR _01314_ VGND net1899 _02957_ sg13g2_o21ai_1
XFILLER_45_439 VPWR VGND sg13g2_decap_8
XFILLER_122_77 VPWR VGND sg13g2_decap_8
X_08699_ VGND VPWR _02911_ net1817 _01337_ _02912_ sg13g2_a21oi_1
X_07719_ _02025_ VPWR _02026_ VGND _01747_ _02024_ sg13g2_o21ai_1
XFILLER_81_770 VPWR VGND sg13g2_decap_8
XFILLER_13_303 VPWR VGND sg13g2_fill_2
X_10730_ _04743_ _04742_ VPWR VGND sg13g2_inv_2
XFILLER_26_697 VPWR VGND sg13g2_fill_2
XFILLER_41_667 VPWR VGND sg13g2_decap_8
XFILLER_40_133 VPWR VGND sg13g2_decap_8
XFILLER_15_42 VPWR VGND sg13g2_decap_8
X_10661_ _04674_ _04670_ _04672_ VPWR VGND sg13g2_nand2_1
XFILLER_25_196 VPWR VGND sg13g2_decap_8
X_12400_ _06242_ _06245_ _06246_ VPWR VGND sg13g2_nor2_1
X_13380_ _07066_ VPWR _00811_ VGND _05367_ _07055_ sg13g2_o21ai_1
XFILLER_12_1009 VPWR VGND sg13g2_decap_4
X_10592_ _04609_ acc_sub.x2\[3\] net1934 VPWR VGND sg13g2_nand2_1
X_12331_ VPWR _06177_ _06176_ VGND sg13g2_inv_1
XFILLER_5_513 VPWR VGND sg13g2_decap_8
XFILLER_126_238 VPWR VGND sg13g2_decap_8
X_12262_ VPWR _06108_ _06078_ VGND sg13g2_inv_1
XFILLER_31_63 VPWR VGND sg13g2_decap_8
XFILLER_108_986 VPWR VGND sg13g2_decap_8
XFILLER_103_0 VPWR VGND sg13g2_decap_8
X_14001_ VPWR _00552_ net87 VGND sg13g2_inv_1
X_11213_ _02959_ _05026_ _05179_ VPWR VGND sg13g2_nor2_1
XFILLER_5_568 VPWR VGND sg13g2_decap_8
X_12193_ _06039_ _06038_ _06027_ VPWR VGND sg13g2_nand2_1
XFILLER_123_967 VPWR VGND sg13g2_decap_8
X_11144_ _05114_ net1698 _05113_ VPWR VGND sg13g2_nand2_1
XFILLER_122_477 VPWR VGND sg13g2_decap_8
XFILLER_110_617 VPWR VGND sg13g2_decap_8
XFILLER_103_680 VPWR VGND sg13g2_decap_8
X_11075_ _04993_ _05046_ _05052_ VPWR VGND sg13g2_nor2_2
XFILLER_48_200 VPWR VGND sg13g2_decap_8
X_14903_ _00704_ VGND VPWR _01423_ acc_sub.op_sign_logic0.mantisa_a\[2\] clknet_5_29__leaf_clk
+ sg13g2_dfrbpq_1
X_10026_ _04114_ _04025_ _04113_ VPWR VGND sg13g2_xnor2_1
XFILLER_76_586 VPWR VGND sg13g2_fill_1
X_14834_ _00635_ VGND VPWR _01358_ state\[0\] clknet_leaf_52_clk sg13g2_dfrbpq_2
XFILLER_17_631 VPWR VGND sg13g2_decap_8
X_14765_ _00566_ VGND VPWR _01289_ acc_sum.exp_mant_logic0.b\[10\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_11977_ _05831_ fpmul.reg_a_out\[10\] fpmul.reg_b_out\[10\] VPWR VGND sg13g2_nand2_1
XFILLER_45_962 VPWR VGND sg13g2_decap_4
X_13716_ VPWR _00267_ net58 VGND sg13g2_inv_1
XFILLER_44_461 VPWR VGND sg13g2_fill_1
X_10928_ net1821 _04933_ _04931_ _04936_ VPWR VGND _04935_ sg13g2_nand4_1
X_14696_ _00497_ VGND VPWR _01224_ fp16_res_pipe.reg_add_sub.q\[0\] clknet_leaf_130_clk
+ sg13g2_dfrbpq_1
X_13647_ VPWR _00198_ net112 VGND sg13g2_inv_1
XFILLER_13_870 VPWR VGND sg13g2_decap_8
X_10859_ VPWR _04871_ _04870_ VGND sg13g2_inv_1
X_13578_ VPWR _00129_ net114 VGND sg13g2_inv_1
X_12529_ _06350_ VPWR _00945_ VGND net1956 _05785_ sg13g2_o21ai_1
XFILLER_9_885 VPWR VGND sg13g2_decap_8
XFILLER_117_238 VPWR VGND sg13g2_decap_8
XFILLER_126_750 VPWR VGND sg13g2_decap_8
XFILLER_114_923 VPWR VGND sg13g2_decap_8
XFILLER_99_623 VPWR VGND sg13g2_fill_2
XFILLER_113_466 VPWR VGND sg13g2_decap_8
XFILLER_99_689 VPWR VGND sg13g2_decap_8
XFILLER_99_667 VPWR VGND sg13g2_fill_1
XFILLER_87_818 VPWR VGND sg13g2_fill_1
XFILLER_101_628 VPWR VGND sg13g2_fill_2
X_09740_ acc_sum.add_renorm0.exp\[3\] _03828_ _03856_ VPWR VGND sg13g2_nor2_1
.ends

